/* -----------------------------------------------------------------------------
 * Part of midgetv
 * 2019. Copyright B. Nossum.
 * For licence, see LICENCE
 * -----------------------------------------------------------------------------ehdr
 * EBR program memory is split into 16-bit wide memory specified here.
 * The memory is up to 4 KiB large
 */
module m_ebr_w16
  # ( parameter EBRAWIDTH = 10,
      parameter [4095:0] prg0 = 4096'h0,
      parameter [4095:0] prg1 = 4096'h0,
      parameter [4095:0] prg2 = 4096'h0,
      parameter [4095:0] prg3 = 4096'h0,
      parameter [4095:0] prg4 = 4096'h0,
      parameter [4095:0] prg5 = 4096'h0,
      parameter [4095:0] prg6 = 4096'h0,
      parameter [4095:0] prg7 = 4096'h0
      )
   (
    input [15:0]          B, //     Output from ALU
    input [EBRAWIDTH-3:0] Rai, //   Read adddress
    input [EBRAWIDTH-3:0] Wai, //   Write adddress
    input                 clk, //   System clock
    input [1:0]           bmask, // Byte masks for write, active LUW
    input                 iwe, //   Write enable
    output [15:0]         DAT_O //  Registered output
    );
   
   localparam NrRamsHere = (1<<(EBRAWIDTH-10));
   
   generate
      
      if ( NrRamsHere == 1 ) begin
         SB_RAM40_4K 
           #(.INIT_0(prg0[ 255:   0]),
             .INIT_1(prg0[ 511: 256]),
             .INIT_2(prg0[ 767: 512]),
             .INIT_3(prg0[1023: 768]),
             .INIT_4(prg0[1279:1024]),
             .INIT_5(prg0[1535:1280]),
             .INIT_6(prg0[1791:1536]),
             .INIT_7(prg0[2047:1792]),
             .INIT_8(prg0[2303:2048]),
             .INIT_9(prg0[2559:2304]),
             .INIT_A(prg0[2815:2560]),
             .INIT_B(prg0[3071:2816]),
             .INIT_C(prg0[3327:3072]),
             .INIT_D(prg0[3583:3328]),
             .INIT_E(prg0[3839:3584]),
             .INIT_F(prg0[4095:3840]))
         mem
           (// Outputs
            .RDATA  ( DAT_O                         ),
            // Input
            .MASK   ( {{8{bmask[1]}},{8{bmask[0]}}} ),
            .WDATA  ( B                             ),
            .WADDR  ( {3'b0,Wai}                    ),
            .RADDR  ( {3'b0,Rai}                    ),
            .RE     ( 1'b1                          ),
            .WE     ( 1'b1                          ),
            .WCLK   ( clk                           ),
            .RCLK   ( clk                           ),
            .RCLKE  ( 1'b1                          ),
            .WCLKE  ( iwe                           )
            /*AUTOINST*/);
         
      end else begin
         /* Split the up to 4 KiB memory into low and high bytes
          */
         localparam [4095:0]
           pb3 = {prg7[4087:4080],prg7[4071:4064],prg7[4055:4048],prg7[4039:4032],prg7[4023:4016],prg7[4007:4000],prg7[3991:3984],prg7[3975:3968],
                  prg7[3959:3952],prg7[3943:3936],prg7[3927:3920],prg7[3911:3904],prg7[3895:3888],prg7[3879:3872],prg7[3863:3856],prg7[3847:3840],
                  prg7[3831:3824],prg7[3815:3808],prg7[3799:3792],prg7[3783:3776],prg7[3767:3760],prg7[3751:3744],prg7[3735:3728],prg7[3719:3712],
                  prg7[3703:3696],prg7[3687:3680],prg7[3671:3664],prg7[3655:3648],prg7[3639:3632],prg7[3623:3616],prg7[3607:3600],prg7[3591:3584],
                  prg7[3575:3568],prg7[3559:3552],prg7[3543:3536],prg7[3527:3520],prg7[3511:3504],prg7[3495:3488],prg7[3479:3472],prg7[3463:3456],
                  prg7[3447:3440],prg7[3431:3424],prg7[3415:3408],prg7[3399:3392],prg7[3383:3376],prg7[3367:3360],prg7[3351:3344],prg7[3335:3328],
                  prg7[3319:3312],prg7[3303:3296],prg7[3287:3280],prg7[3271:3264],prg7[3255:3248],prg7[3239:3232],prg7[3223:3216],prg7[3207:3200],
                  prg7[3191:3184],prg7[3175:3168],prg7[3159:3152],prg7[3143:3136],prg7[3127:3120],prg7[3111:3104],prg7[3095:3088],prg7[3079:3072],
                  prg7[3063:3056],prg7[3047:3040],prg7[3031:3024],prg7[3015:3008],prg7[2999:2992],prg7[2983:2976],prg7[2967:2960],prg7[2951:2944],
                  prg7[2935:2928],prg7[2919:2912],prg7[2903:2896],prg7[2887:2880],prg7[2871:2864],prg7[2855:2848],prg7[2839:2832],prg7[2823:2816],
                  prg7[2807:2800],prg7[2791:2784],prg7[2775:2768],prg7[2759:2752],prg7[2743:2736],prg7[2727:2720],prg7[2711:2704],prg7[2695:2688],
                  prg7[2679:2672],prg7[2663:2656],prg7[2647:2640],prg7[2631:2624],prg7[2615:2608],prg7[2599:2592],prg7[2583:2576],prg7[2567:2560],
                  prg7[2551:2544],prg7[2535:2528],prg7[2519:2512],prg7[2503:2496],prg7[2487:2480],prg7[2471:2464],prg7[2455:2448],prg7[2439:2432],
                  prg7[2423:2416],prg7[2407:2400],prg7[2391:2384],prg7[2375:2368],prg7[2359:2352],prg7[2343:2336],prg7[2327:2320],prg7[2311:2304],
                  prg7[2295:2288],prg7[2279:2272],prg7[2263:2256],prg7[2247:2240],prg7[2231:2224],prg7[2215:2208],prg7[2199:2192],prg7[2183:2176],
                  prg7[2167:2160],prg7[2151:2144],prg7[2135:2128],prg7[2119:2112],prg7[2103:2096],prg7[2087:2080],prg7[2071:2064],prg7[2055:2048],
                  prg7[2039:2032],prg7[2023:2016],prg7[2007:2000],prg7[1991:1984],prg7[1975:1968],prg7[1959:1952],prg7[1943:1936],prg7[1927:1920],
                  prg7[1911:1904],prg7[1895:1888],prg7[1879:1872],prg7[1863:1856],prg7[1847:1840],prg7[1831:1824],prg7[1815:1808],prg7[1799:1792],
                  prg7[1783:1776],prg7[1767:1760],prg7[1751:1744],prg7[1735:1728],prg7[1719:1712],prg7[1703:1696],prg7[1687:1680],prg7[1671:1664],
                  prg7[1655:1648],prg7[1639:1632],prg7[1623:1616],prg7[1607:1600],prg7[1591:1584],prg7[1575:1568],prg7[1559:1552],prg7[1543:1536],
                  prg7[1527:1520],prg7[1511:1504],prg7[1495:1488],prg7[1479:1472],prg7[1463:1456],prg7[1447:1440],prg7[1431:1424],prg7[1415:1408],
                  prg7[1399:1392],prg7[1383:1376],prg7[1367:1360],prg7[1351:1344],prg7[1335:1328],prg7[1319:1312],prg7[1303:1296],prg7[1287:1280],
                  prg7[1271:1264],prg7[1255:1248],prg7[1239:1232],prg7[1223:1216],prg7[1207:1200],prg7[1191:1184],prg7[1175:1168],prg7[1159:1152],
                  prg7[1143:1136],prg7[1127:1120],prg7[1111:1104],prg7[1095:1088],prg7[1079:1072],prg7[1063:1056],prg7[1047:1040],prg7[1031:1024],
                  prg7[1015:1008],prg7[ 999: 992],prg7[ 983: 976],prg7[ 967: 960],prg7[ 951: 944],prg7[ 935: 928],prg7[ 919: 912],prg7[ 903: 896],
                  prg7[ 887: 880],prg7[ 871: 864],prg7[ 855: 848],prg7[ 839: 832],prg7[ 823: 816],prg7[ 807: 800],prg7[ 791: 784],prg7[ 775: 768],
                  prg7[ 759: 752],prg7[ 743: 736],prg7[ 727: 720],prg7[ 711: 704],prg7[ 695: 688],prg7[ 679: 672],prg7[ 663: 656],prg7[ 647: 640],
                  prg7[ 631: 624],prg7[ 615: 608],prg7[ 599: 592],prg7[ 583: 576],prg7[ 567: 560],prg7[ 551: 544],prg7[ 535: 528],prg7[ 519: 512],
                  prg7[ 503: 496],prg7[ 487: 480],prg7[ 471: 464],prg7[ 455: 448],prg7[ 439: 432],prg7[ 423: 416],prg7[ 407: 400],prg7[ 391: 384],
                  prg7[ 375: 368],prg7[ 359: 352],prg7[ 343: 336],prg7[ 327: 320],prg7[ 311: 304],prg7[ 295: 288],prg7[ 279: 272],prg7[ 263: 256],
                  prg7[ 247: 240],prg7[ 231: 224],prg7[ 215: 208],prg7[ 199: 192],prg7[ 183: 176],prg7[ 167: 160],prg7[ 151: 144],prg7[ 135: 128],
                  prg7[ 119: 112],prg7[ 103:  96],prg7[  87:  80],prg7[  71:  64],prg7[  55:  48],prg7[  39:  32],prg7[  23:  16],prg7[   7:   0],
                  prg6[4087:4080],prg6[4071:4064],prg6[4055:4048],prg6[4039:4032],prg6[4023:4016],prg6[4007:4000],prg6[3991:3984],prg6[3975:3968],
                  prg6[3959:3952],prg6[3943:3936],prg6[3927:3920],prg6[3911:3904],prg6[3895:3888],prg6[3879:3872],prg6[3863:3856],prg6[3847:3840],
                  prg6[3831:3824],prg6[3815:3808],prg6[3799:3792],prg6[3783:3776],prg6[3767:3760],prg6[3751:3744],prg6[3735:3728],prg6[3719:3712],
                  prg6[3703:3696],prg6[3687:3680],prg6[3671:3664],prg6[3655:3648],prg6[3639:3632],prg6[3623:3616],prg6[3607:3600],prg6[3591:3584],
                  prg6[3575:3568],prg6[3559:3552],prg6[3543:3536],prg6[3527:3520],prg6[3511:3504],prg6[3495:3488],prg6[3479:3472],prg6[3463:3456],
                  prg6[3447:3440],prg6[3431:3424],prg6[3415:3408],prg6[3399:3392],prg6[3383:3376],prg6[3367:3360],prg6[3351:3344],prg6[3335:3328],
                  prg6[3319:3312],prg6[3303:3296],prg6[3287:3280],prg6[3271:3264],prg6[3255:3248],prg6[3239:3232],prg6[3223:3216],prg6[3207:3200],
                  prg6[3191:3184],prg6[3175:3168],prg6[3159:3152],prg6[3143:3136],prg6[3127:3120],prg6[3111:3104],prg6[3095:3088],prg6[3079:3072],
                  prg6[3063:3056],prg6[3047:3040],prg6[3031:3024],prg6[3015:3008],prg6[2999:2992],prg6[2983:2976],prg6[2967:2960],prg6[2951:2944],
                  prg6[2935:2928],prg6[2919:2912],prg6[2903:2896],prg6[2887:2880],prg6[2871:2864],prg6[2855:2848],prg6[2839:2832],prg6[2823:2816],
                  prg6[2807:2800],prg6[2791:2784],prg6[2775:2768],prg6[2759:2752],prg6[2743:2736],prg6[2727:2720],prg6[2711:2704],prg6[2695:2688],
                  prg6[2679:2672],prg6[2663:2656],prg6[2647:2640],prg6[2631:2624],prg6[2615:2608],prg6[2599:2592],prg6[2583:2576],prg6[2567:2560],
                  prg6[2551:2544],prg6[2535:2528],prg6[2519:2512],prg6[2503:2496],prg6[2487:2480],prg6[2471:2464],prg6[2455:2448],prg6[2439:2432],
                  prg6[2423:2416],prg6[2407:2400],prg6[2391:2384],prg6[2375:2368],prg6[2359:2352],prg6[2343:2336],prg6[2327:2320],prg6[2311:2304],
                  prg6[2295:2288],prg6[2279:2272],prg6[2263:2256],prg6[2247:2240],prg6[2231:2224],prg6[2215:2208],prg6[2199:2192],prg6[2183:2176],
                  prg6[2167:2160],prg6[2151:2144],prg6[2135:2128],prg6[2119:2112],prg6[2103:2096],prg6[2087:2080],prg6[2071:2064],prg6[2055:2048],
                  prg6[2039:2032],prg6[2023:2016],prg6[2007:2000],prg6[1991:1984],prg6[1975:1968],prg6[1959:1952],prg6[1943:1936],prg6[1927:1920],
                  prg6[1911:1904],prg6[1895:1888],prg6[1879:1872],prg6[1863:1856],prg6[1847:1840],prg6[1831:1824],prg6[1815:1808],prg6[1799:1792],
                  prg6[1783:1776],prg6[1767:1760],prg6[1751:1744],prg6[1735:1728],prg6[1719:1712],prg6[1703:1696],prg6[1687:1680],prg6[1671:1664],
                  prg6[1655:1648],prg6[1639:1632],prg6[1623:1616],prg6[1607:1600],prg6[1591:1584],prg6[1575:1568],prg6[1559:1552],prg6[1543:1536],
                  prg6[1527:1520],prg6[1511:1504],prg6[1495:1488],prg6[1479:1472],prg6[1463:1456],prg6[1447:1440],prg6[1431:1424],prg6[1415:1408],
                  prg6[1399:1392],prg6[1383:1376],prg6[1367:1360],prg6[1351:1344],prg6[1335:1328],prg6[1319:1312],prg6[1303:1296],prg6[1287:1280],
                  prg6[1271:1264],prg6[1255:1248],prg6[1239:1232],prg6[1223:1216],prg6[1207:1200],prg6[1191:1184],prg6[1175:1168],prg6[1159:1152],
                  prg6[1143:1136],prg6[1127:1120],prg6[1111:1104],prg6[1095:1088],prg6[1079:1072],prg6[1063:1056],prg6[1047:1040],prg6[1031:1024],
                  prg6[1015:1008],prg6[ 999: 992],prg6[ 983: 976],prg6[ 967: 960],prg6[ 951: 944],prg6[ 935: 928],prg6[ 919: 912],prg6[ 903: 896],
                  prg6[ 887: 880],prg6[ 871: 864],prg6[ 855: 848],prg6[ 839: 832],prg6[ 823: 816],prg6[ 807: 800],prg6[ 791: 784],prg6[ 775: 768],
                  prg6[ 759: 752],prg6[ 743: 736],prg6[ 727: 720],prg6[ 711: 704],prg6[ 695: 688],prg6[ 679: 672],prg6[ 663: 656],prg6[ 647: 640],
                  prg6[ 631: 624],prg6[ 615: 608],prg6[ 599: 592],prg6[ 583: 576],prg6[ 567: 560],prg6[ 551: 544],prg6[ 535: 528],prg6[ 519: 512],
                  prg6[ 503: 496],prg6[ 487: 480],prg6[ 471: 464],prg6[ 455: 448],prg6[ 439: 432],prg6[ 423: 416],prg6[ 407: 400],prg6[ 391: 384],
                  prg6[ 375: 368],prg6[ 359: 352],prg6[ 343: 336],prg6[ 327: 320],prg6[ 311: 304],prg6[ 295: 288],prg6[ 279: 272],prg6[ 263: 256],
                  prg6[ 247: 240],prg6[ 231: 224],prg6[ 215: 208],prg6[ 199: 192],prg6[ 183: 176],prg6[ 167: 160],prg6[ 151: 144],prg6[ 135: 128],
                  prg6[ 119: 112],prg6[ 103:  96],prg6[  87:  80],prg6[  71:  64],prg6[  55:  48],prg6[  39:  32],prg6[  23:  16],prg6[   7:   0]};
         localparam [4095:0]
           pb2 = {prg5[4087:4080],prg5[4071:4064],prg5[4055:4048],prg5[4039:4032],prg5[4023:4016],prg5[4007:4000],prg5[3991:3984],prg5[3975:3968],
                  prg5[3959:3952],prg5[3943:3936],prg5[3927:3920],prg5[3911:3904],prg5[3895:3888],prg5[3879:3872],prg5[3863:3856],prg5[3847:3840],
                  prg5[3831:3824],prg5[3815:3808],prg5[3799:3792],prg5[3783:3776],prg5[3767:3760],prg5[3751:3744],prg5[3735:3728],prg5[3719:3712],
                  prg5[3703:3696],prg5[3687:3680],prg5[3671:3664],prg5[3655:3648],prg5[3639:3632],prg5[3623:3616],prg5[3607:3600],prg5[3591:3584],
                  prg5[3575:3568],prg5[3559:3552],prg5[3543:3536],prg5[3527:3520],prg5[3511:3504],prg5[3495:3488],prg5[3479:3472],prg5[3463:3456],
                  prg5[3447:3440],prg5[3431:3424],prg5[3415:3408],prg5[3399:3392],prg5[3383:3376],prg5[3367:3360],prg5[3351:3344],prg5[3335:3328],
                  prg5[3319:3312],prg5[3303:3296],prg5[3287:3280],prg5[3271:3264],prg5[3255:3248],prg5[3239:3232],prg5[3223:3216],prg5[3207:3200],
                  prg5[3191:3184],prg5[3175:3168],prg5[3159:3152],prg5[3143:3136],prg5[3127:3120],prg5[3111:3104],prg5[3095:3088],prg5[3079:3072],
                  prg5[3063:3056],prg5[3047:3040],prg5[3031:3024],prg5[3015:3008],prg5[2999:2992],prg5[2983:2976],prg5[2967:2960],prg5[2951:2944],
                  prg5[2935:2928],prg5[2919:2912],prg5[2903:2896],prg5[2887:2880],prg5[2871:2864],prg5[2855:2848],prg5[2839:2832],prg5[2823:2816],
                  prg5[2807:2800],prg5[2791:2784],prg5[2775:2768],prg5[2759:2752],prg5[2743:2736],prg5[2727:2720],prg5[2711:2704],prg5[2695:2688],
                  prg5[2679:2672],prg5[2663:2656],prg5[2647:2640],prg5[2631:2624],prg5[2615:2608],prg5[2599:2592],prg5[2583:2576],prg5[2567:2560],
                  prg5[2551:2544],prg5[2535:2528],prg5[2519:2512],prg5[2503:2496],prg5[2487:2480],prg5[2471:2464],prg5[2455:2448],prg5[2439:2432],
                  prg5[2423:2416],prg5[2407:2400],prg5[2391:2384],prg5[2375:2368],prg5[2359:2352],prg5[2343:2336],prg5[2327:2320],prg5[2311:2304],
                  prg5[2295:2288],prg5[2279:2272],prg5[2263:2256],prg5[2247:2240],prg5[2231:2224],prg5[2215:2208],prg5[2199:2192],prg5[2183:2176],
                  prg5[2167:2160],prg5[2151:2144],prg5[2135:2128],prg5[2119:2112],prg5[2103:2096],prg5[2087:2080],prg5[2071:2064],prg5[2055:2048],
                  prg5[2039:2032],prg5[2023:2016],prg5[2007:2000],prg5[1991:1984],prg5[1975:1968],prg5[1959:1952],prg5[1943:1936],prg5[1927:1920],
                  prg5[1911:1904],prg5[1895:1888],prg5[1879:1872],prg5[1863:1856],prg5[1847:1840],prg5[1831:1824],prg5[1815:1808],prg5[1799:1792],
                  prg5[1783:1776],prg5[1767:1760],prg5[1751:1744],prg5[1735:1728],prg5[1719:1712],prg5[1703:1696],prg5[1687:1680],prg5[1671:1664],
                  prg5[1655:1648],prg5[1639:1632],prg5[1623:1616],prg5[1607:1600],prg5[1591:1584],prg5[1575:1568],prg5[1559:1552],prg5[1543:1536],
                  prg5[1527:1520],prg5[1511:1504],prg5[1495:1488],prg5[1479:1472],prg5[1463:1456],prg5[1447:1440],prg5[1431:1424],prg5[1415:1408],
                  prg5[1399:1392],prg5[1383:1376],prg5[1367:1360],prg5[1351:1344],prg5[1335:1328],prg5[1319:1312],prg5[1303:1296],prg5[1287:1280],
                  prg5[1271:1264],prg5[1255:1248],prg5[1239:1232],prg5[1223:1216],prg5[1207:1200],prg5[1191:1184],prg5[1175:1168],prg5[1159:1152],
                  prg5[1143:1136],prg5[1127:1120],prg5[1111:1104],prg5[1095:1088],prg5[1079:1072],prg5[1063:1056],prg5[1047:1040],prg5[1031:1024],
                  prg5[1015:1008],prg5[ 999: 992],prg5[ 983: 976],prg5[ 967: 960],prg5[ 951: 944],prg5[ 935: 928],prg5[ 919: 912],prg5[ 903: 896],
                  prg5[ 887: 880],prg5[ 871: 864],prg5[ 855: 848],prg5[ 839: 832],prg5[ 823: 816],prg5[ 807: 800],prg5[ 791: 784],prg5[ 775: 768],
                  prg5[ 759: 752],prg5[ 743: 736],prg5[ 727: 720],prg5[ 711: 704],prg5[ 695: 688],prg5[ 679: 672],prg5[ 663: 656],prg5[ 647: 640],
                  prg5[ 631: 624],prg5[ 615: 608],prg5[ 599: 592],prg5[ 583: 576],prg5[ 567: 560],prg5[ 551: 544],prg5[ 535: 528],prg5[ 519: 512],
                  prg5[ 503: 496],prg5[ 487: 480],prg5[ 471: 464],prg5[ 455: 448],prg5[ 439: 432],prg5[ 423: 416],prg5[ 407: 400],prg5[ 391: 384],
                  prg5[ 375: 368],prg5[ 359: 352],prg5[ 343: 336],prg5[ 327: 320],prg5[ 311: 304],prg5[ 295: 288],prg5[ 279: 272],prg5[ 263: 256],
                  prg5[ 247: 240],prg5[ 231: 224],prg5[ 215: 208],prg5[ 199: 192],prg5[ 183: 176],prg5[ 167: 160],prg5[ 151: 144],prg5[ 135: 128],
                  prg5[ 119: 112],prg5[ 103:  96],prg5[  87:  80],prg5[  71:  64],prg5[  55:  48],prg5[  39:  32],prg5[  23:  16],prg5[   7:   0],
                  prg4[4087:4080],prg4[4071:4064],prg4[4055:4048],prg4[4039:4032],prg4[4023:4016],prg4[4007:4000],prg4[3991:3984],prg4[3975:3968],
                  prg4[3959:3952],prg4[3943:3936],prg4[3927:3920],prg4[3911:3904],prg4[3895:3888],prg4[3879:3872],prg4[3863:3856],prg4[3847:3840],
                  prg4[3831:3824],prg4[3815:3808],prg4[3799:3792],prg4[3783:3776],prg4[3767:3760],prg4[3751:3744],prg4[3735:3728],prg4[3719:3712],
                  prg4[3703:3696],prg4[3687:3680],prg4[3671:3664],prg4[3655:3648],prg4[3639:3632],prg4[3623:3616],prg4[3607:3600],prg4[3591:3584],
                  prg4[3575:3568],prg4[3559:3552],prg4[3543:3536],prg4[3527:3520],prg4[3511:3504],prg4[3495:3488],prg4[3479:3472],prg4[3463:3456],
                  prg4[3447:3440],prg4[3431:3424],prg4[3415:3408],prg4[3399:3392],prg4[3383:3376],prg4[3367:3360],prg4[3351:3344],prg4[3335:3328],
                  prg4[3319:3312],prg4[3303:3296],prg4[3287:3280],prg4[3271:3264],prg4[3255:3248],prg4[3239:3232],prg4[3223:3216],prg4[3207:3200],
                  prg4[3191:3184],prg4[3175:3168],prg4[3159:3152],prg4[3143:3136],prg4[3127:3120],prg4[3111:3104],prg4[3095:3088],prg4[3079:3072],
                  prg4[3063:3056],prg4[3047:3040],prg4[3031:3024],prg4[3015:3008],prg4[2999:2992],prg4[2983:2976],prg4[2967:2960],prg4[2951:2944],
                  prg4[2935:2928],prg4[2919:2912],prg4[2903:2896],prg4[2887:2880],prg4[2871:2864],prg4[2855:2848],prg4[2839:2832],prg4[2823:2816],
                  prg4[2807:2800],prg4[2791:2784],prg4[2775:2768],prg4[2759:2752],prg4[2743:2736],prg4[2727:2720],prg4[2711:2704],prg4[2695:2688],
                  prg4[2679:2672],prg4[2663:2656],prg4[2647:2640],prg4[2631:2624],prg4[2615:2608],prg4[2599:2592],prg4[2583:2576],prg4[2567:2560],
                  prg4[2551:2544],prg4[2535:2528],prg4[2519:2512],prg4[2503:2496],prg4[2487:2480],prg4[2471:2464],prg4[2455:2448],prg4[2439:2432],
                  prg4[2423:2416],prg4[2407:2400],prg4[2391:2384],prg4[2375:2368],prg4[2359:2352],prg4[2343:2336],prg4[2327:2320],prg4[2311:2304],
                  prg4[2295:2288],prg4[2279:2272],prg4[2263:2256],prg4[2247:2240],prg4[2231:2224],prg4[2215:2208],prg4[2199:2192],prg4[2183:2176],
                  prg4[2167:2160],prg4[2151:2144],prg4[2135:2128],prg4[2119:2112],prg4[2103:2096],prg4[2087:2080],prg4[2071:2064],prg4[2055:2048],
                  prg4[2039:2032],prg4[2023:2016],prg4[2007:2000],prg4[1991:1984],prg4[1975:1968],prg4[1959:1952],prg4[1943:1936],prg4[1927:1920],
                  prg4[1911:1904],prg4[1895:1888],prg4[1879:1872],prg4[1863:1856],prg4[1847:1840],prg4[1831:1824],prg4[1815:1808],prg4[1799:1792],
                  prg4[1783:1776],prg4[1767:1760],prg4[1751:1744],prg4[1735:1728],prg4[1719:1712],prg4[1703:1696],prg4[1687:1680],prg4[1671:1664],
                  prg4[1655:1648],prg4[1639:1632],prg4[1623:1616],prg4[1607:1600],prg4[1591:1584],prg4[1575:1568],prg4[1559:1552],prg4[1543:1536],
                  prg4[1527:1520],prg4[1511:1504],prg4[1495:1488],prg4[1479:1472],prg4[1463:1456],prg4[1447:1440],prg4[1431:1424],prg4[1415:1408],
                  prg4[1399:1392],prg4[1383:1376],prg4[1367:1360],prg4[1351:1344],prg4[1335:1328],prg4[1319:1312],prg4[1303:1296],prg4[1287:1280],
                  prg4[1271:1264],prg4[1255:1248],prg4[1239:1232],prg4[1223:1216],prg4[1207:1200],prg4[1191:1184],prg4[1175:1168],prg4[1159:1152],
                  prg4[1143:1136],prg4[1127:1120],prg4[1111:1104],prg4[1095:1088],prg4[1079:1072],prg4[1063:1056],prg4[1047:1040],prg4[1031:1024],
                  prg4[1015:1008],prg4[ 999: 992],prg4[ 983: 976],prg4[ 967: 960],prg4[ 951: 944],prg4[ 935: 928],prg4[ 919: 912],prg4[ 903: 896],
                  prg4[ 887: 880],prg4[ 871: 864],prg4[ 855: 848],prg4[ 839: 832],prg4[ 823: 816],prg4[ 807: 800],prg4[ 791: 784],prg4[ 775: 768],
                  prg4[ 759: 752],prg4[ 743: 736],prg4[ 727: 720],prg4[ 711: 704],prg4[ 695: 688],prg4[ 679: 672],prg4[ 663: 656],prg4[ 647: 640],
                  prg4[ 631: 624],prg4[ 615: 608],prg4[ 599: 592],prg4[ 583: 576],prg4[ 567: 560],prg4[ 551: 544],prg4[ 535: 528],prg4[ 519: 512],
                  prg4[ 503: 496],prg4[ 487: 480],prg4[ 471: 464],prg4[ 455: 448],prg4[ 439: 432],prg4[ 423: 416],prg4[ 407: 400],prg4[ 391: 384],
                  prg4[ 375: 368],prg4[ 359: 352],prg4[ 343: 336],prg4[ 327: 320],prg4[ 311: 304],prg4[ 295: 288],prg4[ 279: 272],prg4[ 263: 256],
                  prg4[ 247: 240],prg4[ 231: 224],prg4[ 215: 208],prg4[ 199: 192],prg4[ 183: 176],prg4[ 167: 160],prg4[ 151: 144],prg4[ 135: 128],
                  prg4[ 119: 112],prg4[ 103:  96],prg4[  87:  80],prg4[  71:  64],prg4[  55:  48],prg4[  39:  32],prg4[  23:  16],prg4[   7:   0]};
         localparam [4095:0]
           pb1 = {prg3[4087:4080],prg3[4071:4064],prg3[4055:4048],prg3[4039:4032],prg3[4023:4016],prg3[4007:4000],prg3[3991:3984],prg3[3975:3968],
                  prg3[3959:3952],prg3[3943:3936],prg3[3927:3920],prg3[3911:3904],prg3[3895:3888],prg3[3879:3872],prg3[3863:3856],prg3[3847:3840],
                  prg3[3831:3824],prg3[3815:3808],prg3[3799:3792],prg3[3783:3776],prg3[3767:3760],prg3[3751:3744],prg3[3735:3728],prg3[3719:3712],
                  prg3[3703:3696],prg3[3687:3680],prg3[3671:3664],prg3[3655:3648],prg3[3639:3632],prg3[3623:3616],prg3[3607:3600],prg3[3591:3584],
                  prg3[3575:3568],prg3[3559:3552],prg3[3543:3536],prg3[3527:3520],prg3[3511:3504],prg3[3495:3488],prg3[3479:3472],prg3[3463:3456],
                  prg3[3447:3440],prg3[3431:3424],prg3[3415:3408],prg3[3399:3392],prg3[3383:3376],prg3[3367:3360],prg3[3351:3344],prg3[3335:3328],
                  prg3[3319:3312],prg3[3303:3296],prg3[3287:3280],prg3[3271:3264],prg3[3255:3248],prg3[3239:3232],prg3[3223:3216],prg3[3207:3200],
                  prg3[3191:3184],prg3[3175:3168],prg3[3159:3152],prg3[3143:3136],prg3[3127:3120],prg3[3111:3104],prg3[3095:3088],prg3[3079:3072],
                  prg3[3063:3056],prg3[3047:3040],prg3[3031:3024],prg3[3015:3008],prg3[2999:2992],prg3[2983:2976],prg3[2967:2960],prg3[2951:2944],
                  prg3[2935:2928],prg3[2919:2912],prg3[2903:2896],prg3[2887:2880],prg3[2871:2864],prg3[2855:2848],prg3[2839:2832],prg3[2823:2816],
                  prg3[2807:2800],prg3[2791:2784],prg3[2775:2768],prg3[2759:2752],prg3[2743:2736],prg3[2727:2720],prg3[2711:2704],prg3[2695:2688],
                  prg3[2679:2672],prg3[2663:2656],prg3[2647:2640],prg3[2631:2624],prg3[2615:2608],prg3[2599:2592],prg3[2583:2576],prg3[2567:2560],
                  prg3[2551:2544],prg3[2535:2528],prg3[2519:2512],prg3[2503:2496],prg3[2487:2480],prg3[2471:2464],prg3[2455:2448],prg3[2439:2432],
                  prg3[2423:2416],prg3[2407:2400],prg3[2391:2384],prg3[2375:2368],prg3[2359:2352],prg3[2343:2336],prg3[2327:2320],prg3[2311:2304],
                  prg3[2295:2288],prg3[2279:2272],prg3[2263:2256],prg3[2247:2240],prg3[2231:2224],prg3[2215:2208],prg3[2199:2192],prg3[2183:2176],
                  prg3[2167:2160],prg3[2151:2144],prg3[2135:2128],prg3[2119:2112],prg3[2103:2096],prg3[2087:2080],prg3[2071:2064],prg3[2055:2048],
                  prg3[2039:2032],prg3[2023:2016],prg3[2007:2000],prg3[1991:1984],prg3[1975:1968],prg3[1959:1952],prg3[1943:1936],prg3[1927:1920],
                  prg3[1911:1904],prg3[1895:1888],prg3[1879:1872],prg3[1863:1856],prg3[1847:1840],prg3[1831:1824],prg3[1815:1808],prg3[1799:1792],
                  prg3[1783:1776],prg3[1767:1760],prg3[1751:1744],prg3[1735:1728],prg3[1719:1712],prg3[1703:1696],prg3[1687:1680],prg3[1671:1664],
                  prg3[1655:1648],prg3[1639:1632],prg3[1623:1616],prg3[1607:1600],prg3[1591:1584],prg3[1575:1568],prg3[1559:1552],prg3[1543:1536],
                  prg3[1527:1520],prg3[1511:1504],prg3[1495:1488],prg3[1479:1472],prg3[1463:1456],prg3[1447:1440],prg3[1431:1424],prg3[1415:1408],
                  prg3[1399:1392],prg3[1383:1376],prg3[1367:1360],prg3[1351:1344],prg3[1335:1328],prg3[1319:1312],prg3[1303:1296],prg3[1287:1280],
                  prg3[1271:1264],prg3[1255:1248],prg3[1239:1232],prg3[1223:1216],prg3[1207:1200],prg3[1191:1184],prg3[1175:1168],prg3[1159:1152],
                  prg3[1143:1136],prg3[1127:1120],prg3[1111:1104],prg3[1095:1088],prg3[1079:1072],prg3[1063:1056],prg3[1047:1040],prg3[1031:1024],
                  prg3[1015:1008],prg3[ 999: 992],prg3[ 983: 976],prg3[ 967: 960],prg3[ 951: 944],prg3[ 935: 928],prg3[ 919: 912],prg3[ 903: 896],
                  prg3[ 887: 880],prg3[ 871: 864],prg3[ 855: 848],prg3[ 839: 832],prg3[ 823: 816],prg3[ 807: 800],prg3[ 791: 784],prg3[ 775: 768],
                  prg3[ 759: 752],prg3[ 743: 736],prg3[ 727: 720],prg3[ 711: 704],prg3[ 695: 688],prg3[ 679: 672],prg3[ 663: 656],prg3[ 647: 640],
                  prg3[ 631: 624],prg3[ 615: 608],prg3[ 599: 592],prg3[ 583: 576],prg3[ 567: 560],prg3[ 551: 544],prg3[ 535: 528],prg3[ 519: 512],
                  prg3[ 503: 496],prg3[ 487: 480],prg3[ 471: 464],prg3[ 455: 448],prg3[ 439: 432],prg3[ 423: 416],prg3[ 407: 400],prg3[ 391: 384],
                  prg3[ 375: 368],prg3[ 359: 352],prg3[ 343: 336],prg3[ 327: 320],prg3[ 311: 304],prg3[ 295: 288],prg3[ 279: 272],prg3[ 263: 256],
                  prg3[ 247: 240],prg3[ 231: 224],prg3[ 215: 208],prg3[ 199: 192],prg3[ 183: 176],prg3[ 167: 160],prg3[ 151: 144],prg3[ 135: 128],
                  prg3[ 119: 112],prg3[ 103:  96],prg3[  87:  80],prg3[  71:  64],prg3[  55:  48],prg3[  39:  32],prg3[  23:  16],prg3[   7:   0],
                  prg2[4087:4080],prg2[4071:4064],prg2[4055:4048],prg2[4039:4032],prg2[4023:4016],prg2[4007:4000],prg2[3991:3984],prg2[3975:3968],
                  prg2[3959:3952],prg2[3943:3936],prg2[3927:3920],prg2[3911:3904],prg2[3895:3888],prg2[3879:3872],prg2[3863:3856],prg2[3847:3840],
                  prg2[3831:3824],prg2[3815:3808],prg2[3799:3792],prg2[3783:3776],prg2[3767:3760],prg2[3751:3744],prg2[3735:3728],prg2[3719:3712],
                  prg2[3703:3696],prg2[3687:3680],prg2[3671:3664],prg2[3655:3648],prg2[3639:3632],prg2[3623:3616],prg2[3607:3600],prg2[3591:3584],
                  prg2[3575:3568],prg2[3559:3552],prg2[3543:3536],prg2[3527:3520],prg2[3511:3504],prg2[3495:3488],prg2[3479:3472],prg2[3463:3456],
                  prg2[3447:3440],prg2[3431:3424],prg2[3415:3408],prg2[3399:3392],prg2[3383:3376],prg2[3367:3360],prg2[3351:3344],prg2[3335:3328],
                  prg2[3319:3312],prg2[3303:3296],prg2[3287:3280],prg2[3271:3264],prg2[3255:3248],prg2[3239:3232],prg2[3223:3216],prg2[3207:3200],
                  prg2[3191:3184],prg2[3175:3168],prg2[3159:3152],prg2[3143:3136],prg2[3127:3120],prg2[3111:3104],prg2[3095:3088],prg2[3079:3072],
                  prg2[3063:3056],prg2[3047:3040],prg2[3031:3024],prg2[3015:3008],prg2[2999:2992],prg2[2983:2976],prg2[2967:2960],prg2[2951:2944],
                  prg2[2935:2928],prg2[2919:2912],prg2[2903:2896],prg2[2887:2880],prg2[2871:2864],prg2[2855:2848],prg2[2839:2832],prg2[2823:2816],
                  prg2[2807:2800],prg2[2791:2784],prg2[2775:2768],prg2[2759:2752],prg2[2743:2736],prg2[2727:2720],prg2[2711:2704],prg2[2695:2688],
                  prg2[2679:2672],prg2[2663:2656],prg2[2647:2640],prg2[2631:2624],prg2[2615:2608],prg2[2599:2592],prg2[2583:2576],prg2[2567:2560],
                  prg2[2551:2544],prg2[2535:2528],prg2[2519:2512],prg2[2503:2496],prg2[2487:2480],prg2[2471:2464],prg2[2455:2448],prg2[2439:2432],
                  prg2[2423:2416],prg2[2407:2400],prg2[2391:2384],prg2[2375:2368],prg2[2359:2352],prg2[2343:2336],prg2[2327:2320],prg2[2311:2304],
                  prg2[2295:2288],prg2[2279:2272],prg2[2263:2256],prg2[2247:2240],prg2[2231:2224],prg2[2215:2208],prg2[2199:2192],prg2[2183:2176],
                  prg2[2167:2160],prg2[2151:2144],prg2[2135:2128],prg2[2119:2112],prg2[2103:2096],prg2[2087:2080],prg2[2071:2064],prg2[2055:2048],
                  prg2[2039:2032],prg2[2023:2016],prg2[2007:2000],prg2[1991:1984],prg2[1975:1968],prg2[1959:1952],prg2[1943:1936],prg2[1927:1920],
                  prg2[1911:1904],prg2[1895:1888],prg2[1879:1872],prg2[1863:1856],prg2[1847:1840],prg2[1831:1824],prg2[1815:1808],prg2[1799:1792],
                  prg2[1783:1776],prg2[1767:1760],prg2[1751:1744],prg2[1735:1728],prg2[1719:1712],prg2[1703:1696],prg2[1687:1680],prg2[1671:1664],
                  prg2[1655:1648],prg2[1639:1632],prg2[1623:1616],prg2[1607:1600],prg2[1591:1584],prg2[1575:1568],prg2[1559:1552],prg2[1543:1536],
                  prg2[1527:1520],prg2[1511:1504],prg2[1495:1488],prg2[1479:1472],prg2[1463:1456],prg2[1447:1440],prg2[1431:1424],prg2[1415:1408],
                  prg2[1399:1392],prg2[1383:1376],prg2[1367:1360],prg2[1351:1344],prg2[1335:1328],prg2[1319:1312],prg2[1303:1296],prg2[1287:1280],
                  prg2[1271:1264],prg2[1255:1248],prg2[1239:1232],prg2[1223:1216],prg2[1207:1200],prg2[1191:1184],prg2[1175:1168],prg2[1159:1152],
                  prg2[1143:1136],prg2[1127:1120],prg2[1111:1104],prg2[1095:1088],prg2[1079:1072],prg2[1063:1056],prg2[1047:1040],prg2[1031:1024],
                  prg2[1015:1008],prg2[ 999: 992],prg2[ 983: 976],prg2[ 967: 960],prg2[ 951: 944],prg2[ 935: 928],prg2[ 919: 912],prg2[ 903: 896],
                  prg2[ 887: 880],prg2[ 871: 864],prg2[ 855: 848],prg2[ 839: 832],prg2[ 823: 816],prg2[ 807: 800],prg2[ 791: 784],prg2[ 775: 768],
                  prg2[ 759: 752],prg2[ 743: 736],prg2[ 727: 720],prg2[ 711: 704],prg2[ 695: 688],prg2[ 679: 672],prg2[ 663: 656],prg2[ 647: 640],
                  prg2[ 631: 624],prg2[ 615: 608],prg2[ 599: 592],prg2[ 583: 576],prg2[ 567: 560],prg2[ 551: 544],prg2[ 535: 528],prg2[ 519: 512],
                  prg2[ 503: 496],prg2[ 487: 480],prg2[ 471: 464],prg2[ 455: 448],prg2[ 439: 432],prg2[ 423: 416],prg2[ 407: 400],prg2[ 391: 384],
                  prg2[ 375: 368],prg2[ 359: 352],prg2[ 343: 336],prg2[ 327: 320],prg2[ 311: 304],prg2[ 295: 288],prg2[ 279: 272],prg2[ 263: 256],
                  prg2[ 247: 240],prg2[ 231: 224],prg2[ 215: 208],prg2[ 199: 192],prg2[ 183: 176],prg2[ 167: 160],prg2[ 151: 144],prg2[ 135: 128],
                  prg2[ 119: 112],prg2[ 103:  96],prg2[  87:  80],prg2[  71:  64],prg2[  55:  48],prg2[  39:  32],prg2[  23:  16],prg2[   7:   0]};
         localparam [4095:0]
           pb0 = {prg1[4087:4080],prg1[4071:4064],prg1[4055:4048],prg1[4039:4032],prg1[4023:4016],prg1[4007:4000],prg1[3991:3984],prg1[3975:3968],
                  prg1[3959:3952],prg1[3943:3936],prg1[3927:3920],prg1[3911:3904],prg1[3895:3888],prg1[3879:3872],prg1[3863:3856],prg1[3847:3840],
                  prg1[3831:3824],prg1[3815:3808],prg1[3799:3792],prg1[3783:3776],prg1[3767:3760],prg1[3751:3744],prg1[3735:3728],prg1[3719:3712],
                  prg1[3703:3696],prg1[3687:3680],prg1[3671:3664],prg1[3655:3648],prg1[3639:3632],prg1[3623:3616],prg1[3607:3600],prg1[3591:3584],
                  prg1[3575:3568],prg1[3559:3552],prg1[3543:3536],prg1[3527:3520],prg1[3511:3504],prg1[3495:3488],prg1[3479:3472],prg1[3463:3456],
                  prg1[3447:3440],prg1[3431:3424],prg1[3415:3408],prg1[3399:3392],prg1[3383:3376],prg1[3367:3360],prg1[3351:3344],prg1[3335:3328],
                  prg1[3319:3312],prg1[3303:3296],prg1[3287:3280],prg1[3271:3264],prg1[3255:3248],prg1[3239:3232],prg1[3223:3216],prg1[3207:3200],
                  prg1[3191:3184],prg1[3175:3168],prg1[3159:3152],prg1[3143:3136],prg1[3127:3120],prg1[3111:3104],prg1[3095:3088],prg1[3079:3072],
                  prg1[3063:3056],prg1[3047:3040],prg1[3031:3024],prg1[3015:3008],prg1[2999:2992],prg1[2983:2976],prg1[2967:2960],prg1[2951:2944],
                  prg1[2935:2928],prg1[2919:2912],prg1[2903:2896],prg1[2887:2880],prg1[2871:2864],prg1[2855:2848],prg1[2839:2832],prg1[2823:2816],
                  prg1[2807:2800],prg1[2791:2784],prg1[2775:2768],prg1[2759:2752],prg1[2743:2736],prg1[2727:2720],prg1[2711:2704],prg1[2695:2688],
                  prg1[2679:2672],prg1[2663:2656],prg1[2647:2640],prg1[2631:2624],prg1[2615:2608],prg1[2599:2592],prg1[2583:2576],prg1[2567:2560],
                  prg1[2551:2544],prg1[2535:2528],prg1[2519:2512],prg1[2503:2496],prg1[2487:2480],prg1[2471:2464],prg1[2455:2448],prg1[2439:2432],
                  prg1[2423:2416],prg1[2407:2400],prg1[2391:2384],prg1[2375:2368],prg1[2359:2352],prg1[2343:2336],prg1[2327:2320],prg1[2311:2304],
                  prg1[2295:2288],prg1[2279:2272],prg1[2263:2256],prg1[2247:2240],prg1[2231:2224],prg1[2215:2208],prg1[2199:2192],prg1[2183:2176],
                  prg1[2167:2160],prg1[2151:2144],prg1[2135:2128],prg1[2119:2112],prg1[2103:2096],prg1[2087:2080],prg1[2071:2064],prg1[2055:2048],
                  prg1[2039:2032],prg1[2023:2016],prg1[2007:2000],prg1[1991:1984],prg1[1975:1968],prg1[1959:1952],prg1[1943:1936],prg1[1927:1920],
                  prg1[1911:1904],prg1[1895:1888],prg1[1879:1872],prg1[1863:1856],prg1[1847:1840],prg1[1831:1824],prg1[1815:1808],prg1[1799:1792],
                  prg1[1783:1776],prg1[1767:1760],prg1[1751:1744],prg1[1735:1728],prg1[1719:1712],prg1[1703:1696],prg1[1687:1680],prg1[1671:1664],
                  prg1[1655:1648],prg1[1639:1632],prg1[1623:1616],prg1[1607:1600],prg1[1591:1584],prg1[1575:1568],prg1[1559:1552],prg1[1543:1536],
                  prg1[1527:1520],prg1[1511:1504],prg1[1495:1488],prg1[1479:1472],prg1[1463:1456],prg1[1447:1440],prg1[1431:1424],prg1[1415:1408],
                  prg1[1399:1392],prg1[1383:1376],prg1[1367:1360],prg1[1351:1344],prg1[1335:1328],prg1[1319:1312],prg1[1303:1296],prg1[1287:1280],
                  prg1[1271:1264],prg1[1255:1248],prg1[1239:1232],prg1[1223:1216],prg1[1207:1200],prg1[1191:1184],prg1[1175:1168],prg1[1159:1152],
                  prg1[1143:1136],prg1[1127:1120],prg1[1111:1104],prg1[1095:1088],prg1[1079:1072],prg1[1063:1056],prg1[1047:1040],prg1[1031:1024],
                  prg1[1015:1008],prg1[ 999: 992],prg1[ 983: 976],prg1[ 967: 960],prg1[ 951: 944],prg1[ 935: 928],prg1[ 919: 912],prg1[ 903: 896],
                  prg1[ 887: 880],prg1[ 871: 864],prg1[ 855: 848],prg1[ 839: 832],prg1[ 823: 816],prg1[ 807: 800],prg1[ 791: 784],prg1[ 775: 768],
                  prg1[ 759: 752],prg1[ 743: 736],prg1[ 727: 720],prg1[ 711: 704],prg1[ 695: 688],prg1[ 679: 672],prg1[ 663: 656],prg1[ 647: 640],
                  prg1[ 631: 624],prg1[ 615: 608],prg1[ 599: 592],prg1[ 583: 576],prg1[ 567: 560],prg1[ 551: 544],prg1[ 535: 528],prg1[ 519: 512],
                  prg1[ 503: 496],prg1[ 487: 480],prg1[ 471: 464],prg1[ 455: 448],prg1[ 439: 432],prg1[ 423: 416],prg1[ 407: 400],prg1[ 391: 384],
                  prg1[ 375: 368],prg1[ 359: 352],prg1[ 343: 336],prg1[ 327: 320],prg1[ 311: 304],prg1[ 295: 288],prg1[ 279: 272],prg1[ 263: 256],
                  prg1[ 247: 240],prg1[ 231: 224],prg1[ 215: 208],prg1[ 199: 192],prg1[ 183: 176],prg1[ 167: 160],prg1[ 151: 144],prg1[ 135: 128],
                  prg1[ 119: 112],prg1[ 103:  96],prg1[  87:  80],prg1[  71:  64],prg1[  55:  48],prg1[  39:  32],prg1[  23:  16],prg1[   7:   0],
                  prg0[4087:4080],prg0[4071:4064],prg0[4055:4048],prg0[4039:4032],prg0[4023:4016],prg0[4007:4000],prg0[3991:3984],prg0[3975:3968],
                  prg0[3959:3952],prg0[3943:3936],prg0[3927:3920],prg0[3911:3904],prg0[3895:3888],prg0[3879:3872],prg0[3863:3856],prg0[3847:3840],
                  prg0[3831:3824],prg0[3815:3808],prg0[3799:3792],prg0[3783:3776],prg0[3767:3760],prg0[3751:3744],prg0[3735:3728],prg0[3719:3712],
                  prg0[3703:3696],prg0[3687:3680],prg0[3671:3664],prg0[3655:3648],prg0[3639:3632],prg0[3623:3616],prg0[3607:3600],prg0[3591:3584],
                  prg0[3575:3568],prg0[3559:3552],prg0[3543:3536],prg0[3527:3520],prg0[3511:3504],prg0[3495:3488],prg0[3479:3472],prg0[3463:3456],
                  prg0[3447:3440],prg0[3431:3424],prg0[3415:3408],prg0[3399:3392],prg0[3383:3376],prg0[3367:3360],prg0[3351:3344],prg0[3335:3328],
                  prg0[3319:3312],prg0[3303:3296],prg0[3287:3280],prg0[3271:3264],prg0[3255:3248],prg0[3239:3232],prg0[3223:3216],prg0[3207:3200],
                  prg0[3191:3184],prg0[3175:3168],prg0[3159:3152],prg0[3143:3136],prg0[3127:3120],prg0[3111:3104],prg0[3095:3088],prg0[3079:3072],
                  prg0[3063:3056],prg0[3047:3040],prg0[3031:3024],prg0[3015:3008],prg0[2999:2992],prg0[2983:2976],prg0[2967:2960],prg0[2951:2944],
                  prg0[2935:2928],prg0[2919:2912],prg0[2903:2896],prg0[2887:2880],prg0[2871:2864],prg0[2855:2848],prg0[2839:2832],prg0[2823:2816],
                  prg0[2807:2800],prg0[2791:2784],prg0[2775:2768],prg0[2759:2752],prg0[2743:2736],prg0[2727:2720],prg0[2711:2704],prg0[2695:2688],
                  prg0[2679:2672],prg0[2663:2656],prg0[2647:2640],prg0[2631:2624],prg0[2615:2608],prg0[2599:2592],prg0[2583:2576],prg0[2567:2560],
                  prg0[2551:2544],prg0[2535:2528],prg0[2519:2512],prg0[2503:2496],prg0[2487:2480],prg0[2471:2464],prg0[2455:2448],prg0[2439:2432],
                  prg0[2423:2416],prg0[2407:2400],prg0[2391:2384],prg0[2375:2368],prg0[2359:2352],prg0[2343:2336],prg0[2327:2320],prg0[2311:2304],
                  prg0[2295:2288],prg0[2279:2272],prg0[2263:2256],prg0[2247:2240],prg0[2231:2224],prg0[2215:2208],prg0[2199:2192],prg0[2183:2176],
                  prg0[2167:2160],prg0[2151:2144],prg0[2135:2128],prg0[2119:2112],prg0[2103:2096],prg0[2087:2080],prg0[2071:2064],prg0[2055:2048],
                  prg0[2039:2032],prg0[2023:2016],prg0[2007:2000],prg0[1991:1984],prg0[1975:1968],prg0[1959:1952],prg0[1943:1936],prg0[1927:1920],
                  prg0[1911:1904],prg0[1895:1888],prg0[1879:1872],prg0[1863:1856],prg0[1847:1840],prg0[1831:1824],prg0[1815:1808],prg0[1799:1792],
                  prg0[1783:1776],prg0[1767:1760],prg0[1751:1744],prg0[1735:1728],prg0[1719:1712],prg0[1703:1696],prg0[1687:1680],prg0[1671:1664],
                  prg0[1655:1648],prg0[1639:1632],prg0[1623:1616],prg0[1607:1600],prg0[1591:1584],prg0[1575:1568],prg0[1559:1552],prg0[1543:1536],
                  prg0[1527:1520],prg0[1511:1504],prg0[1495:1488],prg0[1479:1472],prg0[1463:1456],prg0[1447:1440],prg0[1431:1424],prg0[1415:1408],
                  prg0[1399:1392],prg0[1383:1376],prg0[1367:1360],prg0[1351:1344],prg0[1335:1328],prg0[1319:1312],prg0[1303:1296],prg0[1287:1280],
                  prg0[1271:1264],prg0[1255:1248],prg0[1239:1232],prg0[1223:1216],prg0[1207:1200],prg0[1191:1184],prg0[1175:1168],prg0[1159:1152],
                  prg0[1143:1136],prg0[1127:1120],prg0[1111:1104],prg0[1095:1088],prg0[1079:1072],prg0[1063:1056],prg0[1047:1040],prg0[1031:1024],
                  prg0[1015:1008],prg0[ 999: 992],prg0[ 983: 976],prg0[ 967: 960],prg0[ 951: 944],prg0[ 935: 928],prg0[ 919: 912],prg0[ 903: 896],
                  prg0[ 887: 880],prg0[ 871: 864],prg0[ 855: 848],prg0[ 839: 832],prg0[ 823: 816],prg0[ 807: 800],prg0[ 791: 784],prg0[ 775: 768],
                  prg0[ 759: 752],prg0[ 743: 736],prg0[ 727: 720],prg0[ 711: 704],prg0[ 695: 688],prg0[ 679: 672],prg0[ 663: 656],prg0[ 647: 640],
                  prg0[ 631: 624],prg0[ 615: 608],prg0[ 599: 592],prg0[ 583: 576],prg0[ 567: 560],prg0[ 551: 544],prg0[ 535: 528],prg0[ 519: 512],
                  prg0[ 503: 496],prg0[ 487: 480],prg0[ 471: 464],prg0[ 455: 448],prg0[ 439: 432],prg0[ 423: 416],prg0[ 407: 400],prg0[ 391: 384],
                  prg0[ 375: 368],prg0[ 359: 352],prg0[ 343: 336],prg0[ 327: 320],prg0[ 311: 304],prg0[ 295: 288],prg0[ 279: 272],prg0[ 263: 256],
                  prg0[ 247: 240],prg0[ 231: 224],prg0[ 215: 208],prg0[ 199: 192],prg0[ 183: 176],prg0[ 167: 160],prg0[ 151: 144],prg0[ 135: 128],
                  prg0[ 119: 112],prg0[ 103:  96],prg0[  87:  80],prg0[  71:  64],prg0[  55:  48],prg0[  39:  32],prg0[  23:  16],prg0[   7:   0]};
         localparam [4095:0]
           ph3 = {prg7[4095:4088],prg7[4079:4072],prg7[4063:4056],prg7[4047:4040],prg7[4031:4024],prg7[4015:4008],prg7[3999:3992],prg7[3983:3976],
                  prg7[3967:3960],prg7[3951:3944],prg7[3935:3928],prg7[3919:3912],prg7[3903:3896],prg7[3887:3880],prg7[3871:3864],prg7[3855:3848],
                  prg7[3839:3832],prg7[3823:3816],prg7[3807:3800],prg7[3791:3784],prg7[3775:3768],prg7[3759:3752],prg7[3743:3736],prg7[3727:3720],
                  prg7[3711:3704],prg7[3695:3688],prg7[3679:3672],prg7[3663:3656],prg7[3647:3640],prg7[3631:3624],prg7[3615:3608],prg7[3599:3592],
                  prg7[3583:3576],prg7[3567:3560],prg7[3551:3544],prg7[3535:3528],prg7[3519:3512],prg7[3503:3496],prg7[3487:3480],prg7[3471:3464],
                  prg7[3455:3448],prg7[3439:3432],prg7[3423:3416],prg7[3407:3400],prg7[3391:3384],prg7[3375:3368],prg7[3359:3352],prg7[3343:3336],
                  prg7[3327:3320],prg7[3311:3304],prg7[3295:3288],prg7[3279:3272],prg7[3263:3256],prg7[3247:3240],prg7[3231:3224],prg7[3215:3208],
                  prg7[3199:3192],prg7[3183:3176],prg7[3167:3160],prg7[3151:3144],prg7[3135:3128],prg7[3119:3112],prg7[3103:3096],prg7[3087:3080],
                  prg7[3071:3064],prg7[3055:3048],prg7[3039:3032],prg7[3023:3016],prg7[3007:3000],prg7[2991:2984],prg7[2975:2968],prg7[2959:2952],
                  prg7[2943:2936],prg7[2927:2920],prg7[2911:2904],prg7[2895:2888],prg7[2879:2872],prg7[2863:2856],prg7[2847:2840],prg7[2831:2824],
                  prg7[2815:2808],prg7[2799:2792],prg7[2783:2776],prg7[2767:2760],prg7[2751:2744],prg7[2735:2728],prg7[2719:2712],prg7[2703:2696],
                  prg7[2687:2680],prg7[2671:2664],prg7[2655:2648],prg7[2639:2632],prg7[2623:2616],prg7[2607:2600],prg7[2591:2584],prg7[2575:2568],
                  prg7[2559:2552],prg7[2543:2536],prg7[2527:2520],prg7[2511:2504],prg7[2495:2488],prg7[2479:2472],prg7[2463:2456],prg7[2447:2440],
                  prg7[2431:2424],prg7[2415:2408],prg7[2399:2392],prg7[2383:2376],prg7[2367:2360],prg7[2351:2344],prg7[2335:2328],prg7[2319:2312],
                  prg7[2303:2296],prg7[2287:2280],prg7[2271:2264],prg7[2255:2248],prg7[2239:2232],prg7[2223:2216],prg7[2207:2200],prg7[2191:2184],
                  prg7[2175:2168],prg7[2159:2152],prg7[2143:2136],prg7[2127:2120],prg7[2111:2104],prg7[2095:2088],prg7[2079:2072],prg7[2063:2056],
                  prg7[2047:2040],prg7[2031:2024],prg7[2015:2008],prg7[1999:1992],prg7[1983:1976],prg7[1967:1960],prg7[1951:1944],prg7[1935:1928],
                  prg7[1919:1912],prg7[1903:1896],prg7[1887:1880],prg7[1871:1864],prg7[1855:1848],prg7[1839:1832],prg7[1823:1816],prg7[1807:1800],
                  prg7[1791:1784],prg7[1775:1768],prg7[1759:1752],prg7[1743:1736],prg7[1727:1720],prg7[1711:1704],prg7[1695:1688],prg7[1679:1672],
                  prg7[1663:1656],prg7[1647:1640],prg7[1631:1624],prg7[1615:1608],prg7[1599:1592],prg7[1583:1576],prg7[1567:1560],prg7[1551:1544],
                  prg7[1535:1528],prg7[1519:1512],prg7[1503:1496],prg7[1487:1480],prg7[1471:1464],prg7[1455:1448],prg7[1439:1432],prg7[1423:1416],
                  prg7[1407:1400],prg7[1391:1384],prg7[1375:1368],prg7[1359:1352],prg7[1343:1336],prg7[1327:1320],prg7[1311:1304],prg7[1295:1288],
                  prg7[1279:1272],prg7[1263:1256],prg7[1247:1240],prg7[1231:1224],prg7[1215:1208],prg7[1199:1192],prg7[1183:1176],prg7[1167:1160],
                  prg7[1151:1144],prg7[1135:1128],prg7[1119:1112],prg7[1103:1096],prg7[1087:1080],prg7[1071:1064],prg7[1055:1048],prg7[1039:1032],
                  prg7[1023:1016],prg7[1007:1000],prg7[ 991: 984],prg7[ 975: 968],prg7[ 959: 952],prg7[ 943: 936],prg7[ 927: 920],prg7[ 911: 904],
                  prg7[ 895: 888],prg7[ 879: 872],prg7[ 863: 856],prg7[ 847: 840],prg7[ 831: 824],prg7[ 815: 808],prg7[ 799: 792],prg7[ 783: 776],
                  prg7[ 767: 760],prg7[ 751: 744],prg7[ 735: 728],prg7[ 719: 712],prg7[ 703: 696],prg7[ 687: 680],prg7[ 671: 664],prg7[ 655: 648],
                  prg7[ 639: 632],prg7[ 623: 616],prg7[ 607: 600],prg7[ 591: 584],prg7[ 575: 568],prg7[ 559: 552],prg7[ 543: 536],prg7[ 527: 520],
                  prg7[ 511: 504],prg7[ 495: 488],prg7[ 479: 472],prg7[ 463: 456],prg7[ 447: 440],prg7[ 431: 424],prg7[ 415: 408],prg7[ 399: 392],
                  prg7[ 383: 376],prg7[ 367: 360],prg7[ 351: 344],prg7[ 335: 328],prg7[ 319: 312],prg7[ 303: 296],prg7[ 287: 280],prg7[ 271: 264],
                  prg7[ 255: 248],prg7[ 239: 232],prg7[ 223: 216],prg7[ 207: 200],prg7[ 191: 184],prg7[ 175: 168],prg7[ 159: 152],prg7[ 143: 136],
                  prg7[ 127: 120],prg7[ 111: 104],prg7[  95:  88],prg7[  79:  72],prg7[  63:  56],prg7[  47:  40],prg7[  31:  24],prg7[  15:   8],
                  prg6[4095:4088],prg6[4079:4072],prg6[4063:4056],prg6[4047:4040],prg6[4031:4024],prg6[4015:4008],prg6[3999:3992],prg6[3983:3976],
                  prg6[3967:3960],prg6[3951:3944],prg6[3935:3928],prg6[3919:3912],prg6[3903:3896],prg6[3887:3880],prg6[3871:3864],prg6[3855:3848],
                  prg6[3839:3832],prg6[3823:3816],prg6[3807:3800],prg6[3791:3784],prg6[3775:3768],prg6[3759:3752],prg6[3743:3736],prg6[3727:3720],
                  prg6[3711:3704],prg6[3695:3688],prg6[3679:3672],prg6[3663:3656],prg6[3647:3640],prg6[3631:3624],prg6[3615:3608],prg6[3599:3592],
                  prg6[3583:3576],prg6[3567:3560],prg6[3551:3544],prg6[3535:3528],prg6[3519:3512],prg6[3503:3496],prg6[3487:3480],prg6[3471:3464],
                  prg6[3455:3448],prg6[3439:3432],prg6[3423:3416],prg6[3407:3400],prg6[3391:3384],prg6[3375:3368],prg6[3359:3352],prg6[3343:3336],
                  prg6[3327:3320],prg6[3311:3304],prg6[3295:3288],prg6[3279:3272],prg6[3263:3256],prg6[3247:3240],prg6[3231:3224],prg6[3215:3208],
                  prg6[3199:3192],prg6[3183:3176],prg6[3167:3160],prg6[3151:3144],prg6[3135:3128],prg6[3119:3112],prg6[3103:3096],prg6[3087:3080],
                  prg6[3071:3064],prg6[3055:3048],prg6[3039:3032],prg6[3023:3016],prg6[3007:3000],prg6[2991:2984],prg6[2975:2968],prg6[2959:2952],
                  prg6[2943:2936],prg6[2927:2920],prg6[2911:2904],prg6[2895:2888],prg6[2879:2872],prg6[2863:2856],prg6[2847:2840],prg6[2831:2824],
                  prg6[2815:2808],prg6[2799:2792],prg6[2783:2776],prg6[2767:2760],prg6[2751:2744],prg6[2735:2728],prg6[2719:2712],prg6[2703:2696],
                  prg6[2687:2680],prg6[2671:2664],prg6[2655:2648],prg6[2639:2632],prg6[2623:2616],prg6[2607:2600],prg6[2591:2584],prg6[2575:2568],
                  prg6[2559:2552],prg6[2543:2536],prg6[2527:2520],prg6[2511:2504],prg6[2495:2488],prg6[2479:2472],prg6[2463:2456],prg6[2447:2440],
                  prg6[2431:2424],prg6[2415:2408],prg6[2399:2392],prg6[2383:2376],prg6[2367:2360],prg6[2351:2344],prg6[2335:2328],prg6[2319:2312],
                  prg6[2303:2296],prg6[2287:2280],prg6[2271:2264],prg6[2255:2248],prg6[2239:2232],prg6[2223:2216],prg6[2207:2200],prg6[2191:2184],
                  prg6[2175:2168],prg6[2159:2152],prg6[2143:2136],prg6[2127:2120],prg6[2111:2104],prg6[2095:2088],prg6[2079:2072],prg6[2063:2056],
                  prg6[2047:2040],prg6[2031:2024],prg6[2015:2008],prg6[1999:1992],prg6[1983:1976],prg6[1967:1960],prg6[1951:1944],prg6[1935:1928],
                  prg6[1919:1912],prg6[1903:1896],prg6[1887:1880],prg6[1871:1864],prg6[1855:1848],prg6[1839:1832],prg6[1823:1816],prg6[1807:1800],
                  prg6[1791:1784],prg6[1775:1768],prg6[1759:1752],prg6[1743:1736],prg6[1727:1720],prg6[1711:1704],prg6[1695:1688],prg6[1679:1672],
                  prg6[1663:1656],prg6[1647:1640],prg6[1631:1624],prg6[1615:1608],prg6[1599:1592],prg6[1583:1576],prg6[1567:1560],prg6[1551:1544],
                  prg6[1535:1528],prg6[1519:1512],prg6[1503:1496],prg6[1487:1480],prg6[1471:1464],prg6[1455:1448],prg6[1439:1432],prg6[1423:1416],
                  prg6[1407:1400],prg6[1391:1384],prg6[1375:1368],prg6[1359:1352],prg6[1343:1336],prg6[1327:1320],prg6[1311:1304],prg6[1295:1288],
                  prg6[1279:1272],prg6[1263:1256],prg6[1247:1240],prg6[1231:1224],prg6[1215:1208],prg6[1199:1192],prg6[1183:1176],prg6[1167:1160],
                  prg6[1151:1144],prg6[1135:1128],prg6[1119:1112],prg6[1103:1096],prg6[1087:1080],prg6[1071:1064],prg6[1055:1048],prg6[1039:1032],
                  prg6[1023:1016],prg6[1007:1000],prg6[ 991: 984],prg6[ 975: 968],prg6[ 959: 952],prg6[ 943: 936],prg6[ 927: 920],prg6[ 911: 904],
                  prg6[ 895: 888],prg6[ 879: 872],prg6[ 863: 856],prg6[ 847: 840],prg6[ 831: 824],prg6[ 815: 808],prg6[ 799: 792],prg6[ 783: 776],
                  prg6[ 767: 760],prg6[ 751: 744],prg6[ 735: 728],prg6[ 719: 712],prg6[ 703: 696],prg6[ 687: 680],prg6[ 671: 664],prg6[ 655: 648],
                  prg6[ 639: 632],prg6[ 623: 616],prg6[ 607: 600],prg6[ 591: 584],prg6[ 575: 568],prg6[ 559: 552],prg6[ 543: 536],prg6[ 527: 520],
                  prg6[ 511: 504],prg6[ 495: 488],prg6[ 479: 472],prg6[ 463: 456],prg6[ 447: 440],prg6[ 431: 424],prg6[ 415: 408],prg6[ 399: 392],
                  prg6[ 383: 376],prg6[ 367: 360],prg6[ 351: 344],prg6[ 335: 328],prg6[ 319: 312],prg6[ 303: 296],prg6[ 287: 280],prg6[ 271: 264],
                  prg6[ 255: 248],prg6[ 239: 232],prg6[ 223: 216],prg6[ 207: 200],prg6[ 191: 184],prg6[ 175: 168],prg6[ 159: 152],prg6[ 143: 136],
                  prg6[ 127: 120],prg6[ 111: 104],prg6[  95:  88],prg6[  79:  72],prg6[  63:  56],prg6[  47:  40],prg6[  31:  24],prg6[  15:   8]};
         localparam [4095:0]
           ph2 = {prg5[4095:4088],prg5[4079:4072],prg5[4063:4056],prg5[4047:4040],prg5[4031:4024],prg5[4015:4008],prg5[3999:3992],prg5[3983:3976],
                  prg5[3967:3960],prg5[3951:3944],prg5[3935:3928],prg5[3919:3912],prg5[3903:3896],prg5[3887:3880],prg5[3871:3864],prg5[3855:3848],
                  prg5[3839:3832],prg5[3823:3816],prg5[3807:3800],prg5[3791:3784],prg5[3775:3768],prg5[3759:3752],prg5[3743:3736],prg5[3727:3720],
                  prg5[3711:3704],prg5[3695:3688],prg5[3679:3672],prg5[3663:3656],prg5[3647:3640],prg5[3631:3624],prg5[3615:3608],prg5[3599:3592],
                  prg5[3583:3576],prg5[3567:3560],prg5[3551:3544],prg5[3535:3528],prg5[3519:3512],prg5[3503:3496],prg5[3487:3480],prg5[3471:3464],
                  prg5[3455:3448],prg5[3439:3432],prg5[3423:3416],prg5[3407:3400],prg5[3391:3384],prg5[3375:3368],prg5[3359:3352],prg5[3343:3336],
                  prg5[3327:3320],prg5[3311:3304],prg5[3295:3288],prg5[3279:3272],prg5[3263:3256],prg5[3247:3240],prg5[3231:3224],prg5[3215:3208],
                  prg5[3199:3192],prg5[3183:3176],prg5[3167:3160],prg5[3151:3144],prg5[3135:3128],prg5[3119:3112],prg5[3103:3096],prg5[3087:3080],
                  prg5[3071:3064],prg5[3055:3048],prg5[3039:3032],prg5[3023:3016],prg5[3007:3000],prg5[2991:2984],prg5[2975:2968],prg5[2959:2952],
                  prg5[2943:2936],prg5[2927:2920],prg5[2911:2904],prg5[2895:2888],prg5[2879:2872],prg5[2863:2856],prg5[2847:2840],prg5[2831:2824],
                  prg5[2815:2808],prg5[2799:2792],prg5[2783:2776],prg5[2767:2760],prg5[2751:2744],prg5[2735:2728],prg5[2719:2712],prg5[2703:2696],
                  prg5[2687:2680],prg5[2671:2664],prg5[2655:2648],prg5[2639:2632],prg5[2623:2616],prg5[2607:2600],prg5[2591:2584],prg5[2575:2568],
                  prg5[2559:2552],prg5[2543:2536],prg5[2527:2520],prg5[2511:2504],prg5[2495:2488],prg5[2479:2472],prg5[2463:2456],prg5[2447:2440],
                  prg5[2431:2424],prg5[2415:2408],prg5[2399:2392],prg5[2383:2376],prg5[2367:2360],prg5[2351:2344],prg5[2335:2328],prg5[2319:2312],
                  prg5[2303:2296],prg5[2287:2280],prg5[2271:2264],prg5[2255:2248],prg5[2239:2232],prg5[2223:2216],prg5[2207:2200],prg5[2191:2184],
                  prg5[2175:2168],prg5[2159:2152],prg5[2143:2136],prg5[2127:2120],prg5[2111:2104],prg5[2095:2088],prg5[2079:2072],prg5[2063:2056],
                  prg5[2047:2040],prg5[2031:2024],prg5[2015:2008],prg5[1999:1992],prg5[1983:1976],prg5[1967:1960],prg5[1951:1944],prg5[1935:1928],
                  prg5[1919:1912],prg5[1903:1896],prg5[1887:1880],prg5[1871:1864],prg5[1855:1848],prg5[1839:1832],prg5[1823:1816],prg5[1807:1800],
                  prg5[1791:1784],prg5[1775:1768],prg5[1759:1752],prg5[1743:1736],prg5[1727:1720],prg5[1711:1704],prg5[1695:1688],prg5[1679:1672],
                  prg5[1663:1656],prg5[1647:1640],prg5[1631:1624],prg5[1615:1608],prg5[1599:1592],prg5[1583:1576],prg5[1567:1560],prg5[1551:1544],
                  prg5[1535:1528],prg5[1519:1512],prg5[1503:1496],prg5[1487:1480],prg5[1471:1464],prg5[1455:1448],prg5[1439:1432],prg5[1423:1416],
                  prg5[1407:1400],prg5[1391:1384],prg5[1375:1368],prg5[1359:1352],prg5[1343:1336],prg5[1327:1320],prg5[1311:1304],prg5[1295:1288],
                  prg5[1279:1272],prg5[1263:1256],prg5[1247:1240],prg5[1231:1224],prg5[1215:1208],prg5[1199:1192],prg5[1183:1176],prg5[1167:1160],
                  prg5[1151:1144],prg5[1135:1128],prg5[1119:1112],prg5[1103:1096],prg5[1087:1080],prg5[1071:1064],prg5[1055:1048],prg5[1039:1032],
                  prg5[1023:1016],prg5[1007:1000],prg5[ 991: 984],prg5[ 975: 968],prg5[ 959: 952],prg5[ 943: 936],prg5[ 927: 920],prg5[ 911: 904],
                  prg5[ 895: 888],prg5[ 879: 872],prg5[ 863: 856],prg5[ 847: 840],prg5[ 831: 824],prg5[ 815: 808],prg5[ 799: 792],prg5[ 783: 776],
                  prg5[ 767: 760],prg5[ 751: 744],prg5[ 735: 728],prg5[ 719: 712],prg5[ 703: 696],prg5[ 687: 680],prg5[ 671: 664],prg5[ 655: 648],
                  prg5[ 639: 632],prg5[ 623: 616],prg5[ 607: 600],prg5[ 591: 584],prg5[ 575: 568],prg5[ 559: 552],prg5[ 543: 536],prg5[ 527: 520],
                  prg5[ 511: 504],prg5[ 495: 488],prg5[ 479: 472],prg5[ 463: 456],prg5[ 447: 440],prg5[ 431: 424],prg5[ 415: 408],prg5[ 399: 392],
                  prg5[ 383: 376],prg5[ 367: 360],prg5[ 351: 344],prg5[ 335: 328],prg5[ 319: 312],prg5[ 303: 296],prg5[ 287: 280],prg5[ 271: 264],
                  prg5[ 255: 248],prg5[ 239: 232],prg5[ 223: 216],prg5[ 207: 200],prg5[ 191: 184],prg5[ 175: 168],prg5[ 159: 152],prg5[ 143: 136],
                  prg5[ 127: 120],prg5[ 111: 104],prg5[  95:  88],prg5[  79:  72],prg5[  63:  56],prg5[  47:  40],prg5[  31:  24],prg5[  15:   8],
                  prg4[4095:4088],prg4[4079:4072],prg4[4063:4056],prg4[4047:4040],prg4[4031:4024],prg4[4015:4008],prg4[3999:3992],prg4[3983:3976],
                  prg4[3967:3960],prg4[3951:3944],prg4[3935:3928],prg4[3919:3912],prg4[3903:3896],prg4[3887:3880],prg4[3871:3864],prg4[3855:3848],
                  prg4[3839:3832],prg4[3823:3816],prg4[3807:3800],prg4[3791:3784],prg4[3775:3768],prg4[3759:3752],prg4[3743:3736],prg4[3727:3720],
                  prg4[3711:3704],prg4[3695:3688],prg4[3679:3672],prg4[3663:3656],prg4[3647:3640],prg4[3631:3624],prg4[3615:3608],prg4[3599:3592],
                  prg4[3583:3576],prg4[3567:3560],prg4[3551:3544],prg4[3535:3528],prg4[3519:3512],prg4[3503:3496],prg4[3487:3480],prg4[3471:3464],
                  prg4[3455:3448],prg4[3439:3432],prg4[3423:3416],prg4[3407:3400],prg4[3391:3384],prg4[3375:3368],prg4[3359:3352],prg4[3343:3336],
                  prg4[3327:3320],prg4[3311:3304],prg4[3295:3288],prg4[3279:3272],prg4[3263:3256],prg4[3247:3240],prg4[3231:3224],prg4[3215:3208],
                  prg4[3199:3192],prg4[3183:3176],prg4[3167:3160],prg4[3151:3144],prg4[3135:3128],prg4[3119:3112],prg4[3103:3096],prg4[3087:3080],
                  prg4[3071:3064],prg4[3055:3048],prg4[3039:3032],prg4[3023:3016],prg4[3007:3000],prg4[2991:2984],prg4[2975:2968],prg4[2959:2952],
                  prg4[2943:2936],prg4[2927:2920],prg4[2911:2904],prg4[2895:2888],prg4[2879:2872],prg4[2863:2856],prg4[2847:2840],prg4[2831:2824],
                  prg4[2815:2808],prg4[2799:2792],prg4[2783:2776],prg4[2767:2760],prg4[2751:2744],prg4[2735:2728],prg4[2719:2712],prg4[2703:2696],
                  prg4[2687:2680],prg4[2671:2664],prg4[2655:2648],prg4[2639:2632],prg4[2623:2616],prg4[2607:2600],prg4[2591:2584],prg4[2575:2568],
                  prg4[2559:2552],prg4[2543:2536],prg4[2527:2520],prg4[2511:2504],prg4[2495:2488],prg4[2479:2472],prg4[2463:2456],prg4[2447:2440],
                  prg4[2431:2424],prg4[2415:2408],prg4[2399:2392],prg4[2383:2376],prg4[2367:2360],prg4[2351:2344],prg4[2335:2328],prg4[2319:2312],
                  prg4[2303:2296],prg4[2287:2280],prg4[2271:2264],prg4[2255:2248],prg4[2239:2232],prg4[2223:2216],prg4[2207:2200],prg4[2191:2184],
                  prg4[2175:2168],prg4[2159:2152],prg4[2143:2136],prg4[2127:2120],prg4[2111:2104],prg4[2095:2088],prg4[2079:2072],prg4[2063:2056],
                  prg4[2047:2040],prg4[2031:2024],prg4[2015:2008],prg4[1999:1992],prg4[1983:1976],prg4[1967:1960],prg4[1951:1944],prg4[1935:1928],
                  prg4[1919:1912],prg4[1903:1896],prg4[1887:1880],prg4[1871:1864],prg4[1855:1848],prg4[1839:1832],prg4[1823:1816],prg4[1807:1800],
                  prg4[1791:1784],prg4[1775:1768],prg4[1759:1752],prg4[1743:1736],prg4[1727:1720],prg4[1711:1704],prg4[1695:1688],prg4[1679:1672],
                  prg4[1663:1656],prg4[1647:1640],prg4[1631:1624],prg4[1615:1608],prg4[1599:1592],prg4[1583:1576],prg4[1567:1560],prg4[1551:1544],
                  prg4[1535:1528],prg4[1519:1512],prg4[1503:1496],prg4[1487:1480],prg4[1471:1464],prg4[1455:1448],prg4[1439:1432],prg4[1423:1416],
                  prg4[1407:1400],prg4[1391:1384],prg4[1375:1368],prg4[1359:1352],prg4[1343:1336],prg4[1327:1320],prg4[1311:1304],prg4[1295:1288],
                  prg4[1279:1272],prg4[1263:1256],prg4[1247:1240],prg4[1231:1224],prg4[1215:1208],prg4[1199:1192],prg4[1183:1176],prg4[1167:1160],
                  prg4[1151:1144],prg4[1135:1128],prg4[1119:1112],prg4[1103:1096],prg4[1087:1080],prg4[1071:1064],prg4[1055:1048],prg4[1039:1032],
                  prg4[1023:1016],prg4[1007:1000],prg4[ 991: 984],prg4[ 975: 968],prg4[ 959: 952],prg4[ 943: 936],prg4[ 927: 920],prg4[ 911: 904],
                  prg4[ 895: 888],prg4[ 879: 872],prg4[ 863: 856],prg4[ 847: 840],prg4[ 831: 824],prg4[ 815: 808],prg4[ 799: 792],prg4[ 783: 776],
                  prg4[ 767: 760],prg4[ 751: 744],prg4[ 735: 728],prg4[ 719: 712],prg4[ 703: 696],prg4[ 687: 680],prg4[ 671: 664],prg4[ 655: 648],
                  prg4[ 639: 632],prg4[ 623: 616],prg4[ 607: 600],prg4[ 591: 584],prg4[ 575: 568],prg4[ 559: 552],prg4[ 543: 536],prg4[ 527: 520],
                  prg4[ 511: 504],prg4[ 495: 488],prg4[ 479: 472],prg4[ 463: 456],prg4[ 447: 440],prg4[ 431: 424],prg4[ 415: 408],prg4[ 399: 392],
                  prg4[ 383: 376],prg4[ 367: 360],prg4[ 351: 344],prg4[ 335: 328],prg4[ 319: 312],prg4[ 303: 296],prg4[ 287: 280],prg4[ 271: 264],
                  prg4[ 255: 248],prg4[ 239: 232],prg4[ 223: 216],prg4[ 207: 200],prg4[ 191: 184],prg4[ 175: 168],prg4[ 159: 152],prg4[ 143: 136],
                  prg4[ 127: 120],prg4[ 111: 104],prg4[  95:  88],prg4[  79:  72],prg4[  63:  56],prg4[  47:  40],prg4[  31:  24],prg4[  15:   8]};
         localparam [4095:0]
           ph1 = {prg3[4095:4088],prg3[4079:4072],prg3[4063:4056],prg3[4047:4040],prg3[4031:4024],prg3[4015:4008],prg3[3999:3992],prg3[3983:3976],
                  prg3[3967:3960],prg3[3951:3944],prg3[3935:3928],prg3[3919:3912],prg3[3903:3896],prg3[3887:3880],prg3[3871:3864],prg3[3855:3848],
                  prg3[3839:3832],prg3[3823:3816],prg3[3807:3800],prg3[3791:3784],prg3[3775:3768],prg3[3759:3752],prg3[3743:3736],prg3[3727:3720],
                  prg3[3711:3704],prg3[3695:3688],prg3[3679:3672],prg3[3663:3656],prg3[3647:3640],prg3[3631:3624],prg3[3615:3608],prg3[3599:3592],
                  prg3[3583:3576],prg3[3567:3560],prg3[3551:3544],prg3[3535:3528],prg3[3519:3512],prg3[3503:3496],prg3[3487:3480],prg3[3471:3464],
                  prg3[3455:3448],prg3[3439:3432],prg3[3423:3416],prg3[3407:3400],prg3[3391:3384],prg3[3375:3368],prg3[3359:3352],prg3[3343:3336],
                  prg3[3327:3320],prg3[3311:3304],prg3[3295:3288],prg3[3279:3272],prg3[3263:3256],prg3[3247:3240],prg3[3231:3224],prg3[3215:3208],
                  prg3[3199:3192],prg3[3183:3176],prg3[3167:3160],prg3[3151:3144],prg3[3135:3128],prg3[3119:3112],prg3[3103:3096],prg3[3087:3080],
                  prg3[3071:3064],prg3[3055:3048],prg3[3039:3032],prg3[3023:3016],prg3[3007:3000],prg3[2991:2984],prg3[2975:2968],prg3[2959:2952],
                  prg3[2943:2936],prg3[2927:2920],prg3[2911:2904],prg3[2895:2888],prg3[2879:2872],prg3[2863:2856],prg3[2847:2840],prg3[2831:2824],
                  prg3[2815:2808],prg3[2799:2792],prg3[2783:2776],prg3[2767:2760],prg3[2751:2744],prg3[2735:2728],prg3[2719:2712],prg3[2703:2696],
                  prg3[2687:2680],prg3[2671:2664],prg3[2655:2648],prg3[2639:2632],prg3[2623:2616],prg3[2607:2600],prg3[2591:2584],prg3[2575:2568],
                  prg3[2559:2552],prg3[2543:2536],prg3[2527:2520],prg3[2511:2504],prg3[2495:2488],prg3[2479:2472],prg3[2463:2456],prg3[2447:2440],
                  prg3[2431:2424],prg3[2415:2408],prg3[2399:2392],prg3[2383:2376],prg3[2367:2360],prg3[2351:2344],prg3[2335:2328],prg3[2319:2312],
                  prg3[2303:2296],prg3[2287:2280],prg3[2271:2264],prg3[2255:2248],prg3[2239:2232],prg3[2223:2216],prg3[2207:2200],prg3[2191:2184],
                  prg3[2175:2168],prg3[2159:2152],prg3[2143:2136],prg3[2127:2120],prg3[2111:2104],prg3[2095:2088],prg3[2079:2072],prg3[2063:2056],
                  prg3[2047:2040],prg3[2031:2024],prg3[2015:2008],prg3[1999:1992],prg3[1983:1976],prg3[1967:1960],prg3[1951:1944],prg3[1935:1928],
                  prg3[1919:1912],prg3[1903:1896],prg3[1887:1880],prg3[1871:1864],prg3[1855:1848],prg3[1839:1832],prg3[1823:1816],prg3[1807:1800],
                  prg3[1791:1784],prg3[1775:1768],prg3[1759:1752],prg3[1743:1736],prg3[1727:1720],prg3[1711:1704],prg3[1695:1688],prg3[1679:1672],
                  prg3[1663:1656],prg3[1647:1640],prg3[1631:1624],prg3[1615:1608],prg3[1599:1592],prg3[1583:1576],prg3[1567:1560],prg3[1551:1544],
                  prg3[1535:1528],prg3[1519:1512],prg3[1503:1496],prg3[1487:1480],prg3[1471:1464],prg3[1455:1448],prg3[1439:1432],prg3[1423:1416],
                  prg3[1407:1400],prg3[1391:1384],prg3[1375:1368],prg3[1359:1352],prg3[1343:1336],prg3[1327:1320],prg3[1311:1304],prg3[1295:1288],
                  prg3[1279:1272],prg3[1263:1256],prg3[1247:1240],prg3[1231:1224],prg3[1215:1208],prg3[1199:1192],prg3[1183:1176],prg3[1167:1160],
                  prg3[1151:1144],prg3[1135:1128],prg3[1119:1112],prg3[1103:1096],prg3[1087:1080],prg3[1071:1064],prg3[1055:1048],prg3[1039:1032],
                  prg3[1023:1016],prg3[1007:1000],prg3[ 991: 984],prg3[ 975: 968],prg3[ 959: 952],prg3[ 943: 936],prg3[ 927: 920],prg3[ 911: 904],
                  prg3[ 895: 888],prg3[ 879: 872],prg3[ 863: 856],prg3[ 847: 840],prg3[ 831: 824],prg3[ 815: 808],prg3[ 799: 792],prg3[ 783: 776],
                  prg3[ 767: 760],prg3[ 751: 744],prg3[ 735: 728],prg3[ 719: 712],prg3[ 703: 696],prg3[ 687: 680],prg3[ 671: 664],prg3[ 655: 648],
                  prg3[ 639: 632],prg3[ 623: 616],prg3[ 607: 600],prg3[ 591: 584],prg3[ 575: 568],prg3[ 559: 552],prg3[ 543: 536],prg3[ 527: 520],
                  prg3[ 511: 504],prg3[ 495: 488],prg3[ 479: 472],prg3[ 463: 456],prg3[ 447: 440],prg3[ 431: 424],prg3[ 415: 408],prg3[ 399: 392],
                  prg3[ 383: 376],prg3[ 367: 360],prg3[ 351: 344],prg3[ 335: 328],prg3[ 319: 312],prg3[ 303: 296],prg3[ 287: 280],prg3[ 271: 264],
                  prg3[ 255: 248],prg3[ 239: 232],prg3[ 223: 216],prg3[ 207: 200],prg3[ 191: 184],prg3[ 175: 168],prg3[ 159: 152],prg3[ 143: 136],
                  prg3[ 127: 120],prg3[ 111: 104],prg3[  95:  88],prg3[  79:  72],prg3[  63:  56],prg3[  47:  40],prg3[  31:  24],prg3[  15:   8],
                  prg2[4095:4088],prg2[4079:4072],prg2[4063:4056],prg2[4047:4040],prg2[4031:4024],prg2[4015:4008],prg2[3999:3992],prg2[3983:3976],
                  prg2[3967:3960],prg2[3951:3944],prg2[3935:3928],prg2[3919:3912],prg2[3903:3896],prg2[3887:3880],prg2[3871:3864],prg2[3855:3848],
                  prg2[3839:3832],prg2[3823:3816],prg2[3807:3800],prg2[3791:3784],prg2[3775:3768],prg2[3759:3752],prg2[3743:3736],prg2[3727:3720],
                  prg2[3711:3704],prg2[3695:3688],prg2[3679:3672],prg2[3663:3656],prg2[3647:3640],prg2[3631:3624],prg2[3615:3608],prg2[3599:3592],
                  prg2[3583:3576],prg2[3567:3560],prg2[3551:3544],prg2[3535:3528],prg2[3519:3512],prg2[3503:3496],prg2[3487:3480],prg2[3471:3464],
                  prg2[3455:3448],prg2[3439:3432],prg2[3423:3416],prg2[3407:3400],prg2[3391:3384],prg2[3375:3368],prg2[3359:3352],prg2[3343:3336],
                  prg2[3327:3320],prg2[3311:3304],prg2[3295:3288],prg2[3279:3272],prg2[3263:3256],prg2[3247:3240],prg2[3231:3224],prg2[3215:3208],
                  prg2[3199:3192],prg2[3183:3176],prg2[3167:3160],prg2[3151:3144],prg2[3135:3128],prg2[3119:3112],prg2[3103:3096],prg2[3087:3080],
                  prg2[3071:3064],prg2[3055:3048],prg2[3039:3032],prg2[3023:3016],prg2[3007:3000],prg2[2991:2984],prg2[2975:2968],prg2[2959:2952],
                  prg2[2943:2936],prg2[2927:2920],prg2[2911:2904],prg2[2895:2888],prg2[2879:2872],prg2[2863:2856],prg2[2847:2840],prg2[2831:2824],
                  prg2[2815:2808],prg2[2799:2792],prg2[2783:2776],prg2[2767:2760],prg2[2751:2744],prg2[2735:2728],prg2[2719:2712],prg2[2703:2696],
                  prg2[2687:2680],prg2[2671:2664],prg2[2655:2648],prg2[2639:2632],prg2[2623:2616],prg2[2607:2600],prg2[2591:2584],prg2[2575:2568],
                  prg2[2559:2552],prg2[2543:2536],prg2[2527:2520],prg2[2511:2504],prg2[2495:2488],prg2[2479:2472],prg2[2463:2456],prg2[2447:2440],
                  prg2[2431:2424],prg2[2415:2408],prg2[2399:2392],prg2[2383:2376],prg2[2367:2360],prg2[2351:2344],prg2[2335:2328],prg2[2319:2312],
                  prg2[2303:2296],prg2[2287:2280],prg2[2271:2264],prg2[2255:2248],prg2[2239:2232],prg2[2223:2216],prg2[2207:2200],prg2[2191:2184],
                  prg2[2175:2168],prg2[2159:2152],prg2[2143:2136],prg2[2127:2120],prg2[2111:2104],prg2[2095:2088],prg2[2079:2072],prg2[2063:2056],
                  prg2[2047:2040],prg2[2031:2024],prg2[2015:2008],prg2[1999:1992],prg2[1983:1976],prg2[1967:1960],prg2[1951:1944],prg2[1935:1928],
                  prg2[1919:1912],prg2[1903:1896],prg2[1887:1880],prg2[1871:1864],prg2[1855:1848],prg2[1839:1832],prg2[1823:1816],prg2[1807:1800],
                  prg2[1791:1784],prg2[1775:1768],prg2[1759:1752],prg2[1743:1736],prg2[1727:1720],prg2[1711:1704],prg2[1695:1688],prg2[1679:1672],
                  prg2[1663:1656],prg2[1647:1640],prg2[1631:1624],prg2[1615:1608],prg2[1599:1592],prg2[1583:1576],prg2[1567:1560],prg2[1551:1544],
                  prg2[1535:1528],prg2[1519:1512],prg2[1503:1496],prg2[1487:1480],prg2[1471:1464],prg2[1455:1448],prg2[1439:1432],prg2[1423:1416],
                  prg2[1407:1400],prg2[1391:1384],prg2[1375:1368],prg2[1359:1352],prg2[1343:1336],prg2[1327:1320],prg2[1311:1304],prg2[1295:1288],
                  prg2[1279:1272],prg2[1263:1256],prg2[1247:1240],prg2[1231:1224],prg2[1215:1208],prg2[1199:1192],prg2[1183:1176],prg2[1167:1160],
                  prg2[1151:1144],prg2[1135:1128],prg2[1119:1112],prg2[1103:1096],prg2[1087:1080],prg2[1071:1064],prg2[1055:1048],prg2[1039:1032],
                  prg2[1023:1016],prg2[1007:1000],prg2[ 991: 984],prg2[ 975: 968],prg2[ 959: 952],prg2[ 943: 936],prg2[ 927: 920],prg2[ 911: 904],
                  prg2[ 895: 888],prg2[ 879: 872],prg2[ 863: 856],prg2[ 847: 840],prg2[ 831: 824],prg2[ 815: 808],prg2[ 799: 792],prg2[ 783: 776],
                  prg2[ 767: 760],prg2[ 751: 744],prg2[ 735: 728],prg2[ 719: 712],prg2[ 703: 696],prg2[ 687: 680],prg2[ 671: 664],prg2[ 655: 648],
                  prg2[ 639: 632],prg2[ 623: 616],prg2[ 607: 600],prg2[ 591: 584],prg2[ 575: 568],prg2[ 559: 552],prg2[ 543: 536],prg2[ 527: 520],
                  prg2[ 511: 504],prg2[ 495: 488],prg2[ 479: 472],prg2[ 463: 456],prg2[ 447: 440],prg2[ 431: 424],prg2[ 415: 408],prg2[ 399: 392],
                  prg2[ 383: 376],prg2[ 367: 360],prg2[ 351: 344],prg2[ 335: 328],prg2[ 319: 312],prg2[ 303: 296],prg2[ 287: 280],prg2[ 271: 264],
                  prg2[ 255: 248],prg2[ 239: 232],prg2[ 223: 216],prg2[ 207: 200],prg2[ 191: 184],prg2[ 175: 168],prg2[ 159: 152],prg2[ 143: 136],
                  prg2[ 127: 120],prg2[ 111: 104],prg2[  95:  88],prg2[  79:  72],prg2[  63:  56],prg2[  47:  40],prg2[  31:  24],prg2[  15:   8]};
         localparam [4095:0]
           ph0 = {prg1[4095:4088],prg1[4079:4072],prg1[4063:4056],prg1[4047:4040],prg1[4031:4024],prg1[4015:4008],prg1[3999:3992],prg1[3983:3976],
                  prg1[3967:3960],prg1[3951:3944],prg1[3935:3928],prg1[3919:3912],prg1[3903:3896],prg1[3887:3880],prg1[3871:3864],prg1[3855:3848],
                  prg1[3839:3832],prg1[3823:3816],prg1[3807:3800],prg1[3791:3784],prg1[3775:3768],prg1[3759:3752],prg1[3743:3736],prg1[3727:3720],
                  prg1[3711:3704],prg1[3695:3688],prg1[3679:3672],prg1[3663:3656],prg1[3647:3640],prg1[3631:3624],prg1[3615:3608],prg1[3599:3592],
                  prg1[3583:3576],prg1[3567:3560],prg1[3551:3544],prg1[3535:3528],prg1[3519:3512],prg1[3503:3496],prg1[3487:3480],prg1[3471:3464],
                  prg1[3455:3448],prg1[3439:3432],prg1[3423:3416],prg1[3407:3400],prg1[3391:3384],prg1[3375:3368],prg1[3359:3352],prg1[3343:3336],
                  prg1[3327:3320],prg1[3311:3304],prg1[3295:3288],prg1[3279:3272],prg1[3263:3256],prg1[3247:3240],prg1[3231:3224],prg1[3215:3208],
                  prg1[3199:3192],prg1[3183:3176],prg1[3167:3160],prg1[3151:3144],prg1[3135:3128],prg1[3119:3112],prg1[3103:3096],prg1[3087:3080],
                  prg1[3071:3064],prg1[3055:3048],prg1[3039:3032],prg1[3023:3016],prg1[3007:3000],prg1[2991:2984],prg1[2975:2968],prg1[2959:2952],
                  prg1[2943:2936],prg1[2927:2920],prg1[2911:2904],prg1[2895:2888],prg1[2879:2872],prg1[2863:2856],prg1[2847:2840],prg1[2831:2824],
                  prg1[2815:2808],prg1[2799:2792],prg1[2783:2776],prg1[2767:2760],prg1[2751:2744],prg1[2735:2728],prg1[2719:2712],prg1[2703:2696],
                  prg1[2687:2680],prg1[2671:2664],prg1[2655:2648],prg1[2639:2632],prg1[2623:2616],prg1[2607:2600],prg1[2591:2584],prg1[2575:2568],
                  prg1[2559:2552],prg1[2543:2536],prg1[2527:2520],prg1[2511:2504],prg1[2495:2488],prg1[2479:2472],prg1[2463:2456],prg1[2447:2440],
                  prg1[2431:2424],prg1[2415:2408],prg1[2399:2392],prg1[2383:2376],prg1[2367:2360],prg1[2351:2344],prg1[2335:2328],prg1[2319:2312],
                  prg1[2303:2296],prg1[2287:2280],prg1[2271:2264],prg1[2255:2248],prg1[2239:2232],prg1[2223:2216],prg1[2207:2200],prg1[2191:2184],
                  prg1[2175:2168],prg1[2159:2152],prg1[2143:2136],prg1[2127:2120],prg1[2111:2104],prg1[2095:2088],prg1[2079:2072],prg1[2063:2056],
                  prg1[2047:2040],prg1[2031:2024],prg1[2015:2008],prg1[1999:1992],prg1[1983:1976],prg1[1967:1960],prg1[1951:1944],prg1[1935:1928],
                  prg1[1919:1912],prg1[1903:1896],prg1[1887:1880],prg1[1871:1864],prg1[1855:1848],prg1[1839:1832],prg1[1823:1816],prg1[1807:1800],
                  prg1[1791:1784],prg1[1775:1768],prg1[1759:1752],prg1[1743:1736],prg1[1727:1720],prg1[1711:1704],prg1[1695:1688],prg1[1679:1672],
                  prg1[1663:1656],prg1[1647:1640],prg1[1631:1624],prg1[1615:1608],prg1[1599:1592],prg1[1583:1576],prg1[1567:1560],prg1[1551:1544],
                  prg1[1535:1528],prg1[1519:1512],prg1[1503:1496],prg1[1487:1480],prg1[1471:1464],prg1[1455:1448],prg1[1439:1432],prg1[1423:1416],
                  prg1[1407:1400],prg1[1391:1384],prg1[1375:1368],prg1[1359:1352],prg1[1343:1336],prg1[1327:1320],prg1[1311:1304],prg1[1295:1288],
                  prg1[1279:1272],prg1[1263:1256],prg1[1247:1240],prg1[1231:1224],prg1[1215:1208],prg1[1199:1192],prg1[1183:1176],prg1[1167:1160],
                  prg1[1151:1144],prg1[1135:1128],prg1[1119:1112],prg1[1103:1096],prg1[1087:1080],prg1[1071:1064],prg1[1055:1048],prg1[1039:1032],
                  prg1[1023:1016],prg1[1007:1000],prg1[ 991: 984],prg1[ 975: 968],prg1[ 959: 952],prg1[ 943: 936],prg1[ 927: 920],prg1[ 911: 904],
                  prg1[ 895: 888],prg1[ 879: 872],prg1[ 863: 856],prg1[ 847: 840],prg1[ 831: 824],prg1[ 815: 808],prg1[ 799: 792],prg1[ 783: 776],
                  prg1[ 767: 760],prg1[ 751: 744],prg1[ 735: 728],prg1[ 719: 712],prg1[ 703: 696],prg1[ 687: 680],prg1[ 671: 664],prg1[ 655: 648],
                  prg1[ 639: 632],prg1[ 623: 616],prg1[ 607: 600],prg1[ 591: 584],prg1[ 575: 568],prg1[ 559: 552],prg1[ 543: 536],prg1[ 527: 520],
                  prg1[ 511: 504],prg1[ 495: 488],prg1[ 479: 472],prg1[ 463: 456],prg1[ 447: 440],prg1[ 431: 424],prg1[ 415: 408],prg1[ 399: 392],
                  prg1[ 383: 376],prg1[ 367: 360],prg1[ 351: 344],prg1[ 335: 328],prg1[ 319: 312],prg1[ 303: 296],prg1[ 287: 280],prg1[ 271: 264],
                  prg1[ 255: 248],prg1[ 239: 232],prg1[ 223: 216],prg1[ 207: 200],prg1[ 191: 184],prg1[ 175: 168],prg1[ 159: 152],prg1[ 143: 136],
                  prg1[ 127: 120],prg1[ 111: 104],prg1[  95:  88],prg1[  79:  72],prg1[  63:  56],prg1[  47:  40],prg1[  31:  24],prg1[  15:   8],
                  prg0[4095:4088],prg0[4079:4072],prg0[4063:4056],prg0[4047:4040],prg0[4031:4024],prg0[4015:4008],prg0[3999:3992],prg0[3983:3976],
                  prg0[3967:3960],prg0[3951:3944],prg0[3935:3928],prg0[3919:3912],prg0[3903:3896],prg0[3887:3880],prg0[3871:3864],prg0[3855:3848],
                  prg0[3839:3832],prg0[3823:3816],prg0[3807:3800],prg0[3791:3784],prg0[3775:3768],prg0[3759:3752],prg0[3743:3736],prg0[3727:3720],
                  prg0[3711:3704],prg0[3695:3688],prg0[3679:3672],prg0[3663:3656],prg0[3647:3640],prg0[3631:3624],prg0[3615:3608],prg0[3599:3592],
                  prg0[3583:3576],prg0[3567:3560],prg0[3551:3544],prg0[3535:3528],prg0[3519:3512],prg0[3503:3496],prg0[3487:3480],prg0[3471:3464],
                  prg0[3455:3448],prg0[3439:3432],prg0[3423:3416],prg0[3407:3400],prg0[3391:3384],prg0[3375:3368],prg0[3359:3352],prg0[3343:3336],
                  prg0[3327:3320],prg0[3311:3304],prg0[3295:3288],prg0[3279:3272],prg0[3263:3256],prg0[3247:3240],prg0[3231:3224],prg0[3215:3208],
                  prg0[3199:3192],prg0[3183:3176],prg0[3167:3160],prg0[3151:3144],prg0[3135:3128],prg0[3119:3112],prg0[3103:3096],prg0[3087:3080],
                  prg0[3071:3064],prg0[3055:3048],prg0[3039:3032],prg0[3023:3016],prg0[3007:3000],prg0[2991:2984],prg0[2975:2968],prg0[2959:2952],
                  prg0[2943:2936],prg0[2927:2920],prg0[2911:2904],prg0[2895:2888],prg0[2879:2872],prg0[2863:2856],prg0[2847:2840],prg0[2831:2824],
                  prg0[2815:2808],prg0[2799:2792],prg0[2783:2776],prg0[2767:2760],prg0[2751:2744],prg0[2735:2728],prg0[2719:2712],prg0[2703:2696],
                  prg0[2687:2680],prg0[2671:2664],prg0[2655:2648],prg0[2639:2632],prg0[2623:2616],prg0[2607:2600],prg0[2591:2584],prg0[2575:2568],
                  prg0[2559:2552],prg0[2543:2536],prg0[2527:2520],prg0[2511:2504],prg0[2495:2488],prg0[2479:2472],prg0[2463:2456],prg0[2447:2440],
                  prg0[2431:2424],prg0[2415:2408],prg0[2399:2392],prg0[2383:2376],prg0[2367:2360],prg0[2351:2344],prg0[2335:2328],prg0[2319:2312],
                  prg0[2303:2296],prg0[2287:2280],prg0[2271:2264],prg0[2255:2248],prg0[2239:2232],prg0[2223:2216],prg0[2207:2200],prg0[2191:2184],
                  prg0[2175:2168],prg0[2159:2152],prg0[2143:2136],prg0[2127:2120],prg0[2111:2104],prg0[2095:2088],prg0[2079:2072],prg0[2063:2056],
                  prg0[2047:2040],prg0[2031:2024],prg0[2015:2008],prg0[1999:1992],prg0[1983:1976],prg0[1967:1960],prg0[1951:1944],prg0[1935:1928],
                  prg0[1919:1912],prg0[1903:1896],prg0[1887:1880],prg0[1871:1864],prg0[1855:1848],prg0[1839:1832],prg0[1823:1816],prg0[1807:1800],
                  prg0[1791:1784],prg0[1775:1768],prg0[1759:1752],prg0[1743:1736],prg0[1727:1720],prg0[1711:1704],prg0[1695:1688],prg0[1679:1672],
                  prg0[1663:1656],prg0[1647:1640],prg0[1631:1624],prg0[1615:1608],prg0[1599:1592],prg0[1583:1576],prg0[1567:1560],prg0[1551:1544],
                  prg0[1535:1528],prg0[1519:1512],prg0[1503:1496],prg0[1487:1480],prg0[1471:1464],prg0[1455:1448],prg0[1439:1432],prg0[1423:1416],
                  prg0[1407:1400],prg0[1391:1384],prg0[1375:1368],prg0[1359:1352],prg0[1343:1336],prg0[1327:1320],prg0[1311:1304],prg0[1295:1288],
                  prg0[1279:1272],prg0[1263:1256],prg0[1247:1240],prg0[1231:1224],prg0[1215:1208],prg0[1199:1192],prg0[1183:1176],prg0[1167:1160],
                  prg0[1151:1144],prg0[1135:1128],prg0[1119:1112],prg0[1103:1096],prg0[1087:1080],prg0[1071:1064],prg0[1055:1048],prg0[1039:1032],
                  prg0[1023:1016],prg0[1007:1000],prg0[ 991: 984],prg0[ 975: 968],prg0[ 959: 952],prg0[ 943: 936],prg0[ 927: 920],prg0[ 911: 904],
                  prg0[ 895: 888],prg0[ 879: 872],prg0[ 863: 856],prg0[ 847: 840],prg0[ 831: 824],prg0[ 815: 808],prg0[ 799: 792],prg0[ 783: 776],
                  prg0[ 767: 760],prg0[ 751: 744],prg0[ 735: 728],prg0[ 719: 712],prg0[ 703: 696],prg0[ 687: 680],prg0[ 671: 664],prg0[ 655: 648],
                  prg0[ 639: 632],prg0[ 623: 616],prg0[ 607: 600],prg0[ 591: 584],prg0[ 575: 568],prg0[ 559: 552],prg0[ 543: 536],prg0[ 527: 520],
                  prg0[ 511: 504],prg0[ 495: 488],prg0[ 479: 472],prg0[ 463: 456],prg0[ 447: 440],prg0[ 431: 424],prg0[ 415: 408],prg0[ 399: 392],
                  prg0[ 383: 376],prg0[ 367: 360],prg0[ 351: 344],prg0[ 335: 328],prg0[ 319: 312],prg0[ 303: 296],prg0[ 287: 280],prg0[ 271: 264],
                  prg0[ 255: 248],prg0[ 239: 232],prg0[ 223: 216],prg0[ 207: 200],prg0[ 191: 184],prg0[ 175: 168],prg0[ 159: 152],prg0[ 143: 136],
                  prg0[ 127: 120],prg0[ 111: 104],prg0[  95:  88],prg0[  79:  72],prg0[  63:  56],prg0[  47:  40],prg0[  31:  24],prg0[  15:   8]};

         m_ebr_w8 #(.EBRAWIDTH(EBRAWIDTH),
                    .prg0(pb0), .prg1(pb1), .prg2(pb2), .prg3(pb3))
         ebrb 
           (// Inputs
            .bmask                      (bmask[0]),
            /*AUTOINST*/
            // Outputs
            .DAT_O                      (DAT_O[7:0]),
            // Inputs
            .B                          (B[7:0]),
            .Rai                        (Rai[EBRAWIDTH-3:0]),
            .Wai                        (Wai[EBRAWIDTH-3:0]),
            .clk                        (clk),
            .iwe                        (iwe));
   
         m_ebr_w8 #(.EBRAWIDTH(EBRAWIDTH),
                    .prg0(ph0), .prg1(ph1), .prg2(ph2), .prg3(ph3))
         ebrh
           (// Outputs
            .DAT_O                      (DAT_O[15:8]),
            // Inputs
            .B                          (B[15:8]),
            .bmask                      (bmask[1]),
            /*AUTOINST*/
            // Inputs
            .Rai                        (Rai[EBRAWIDTH-3:0]),
            .Wai                        (Wai[EBRAWIDTH-3:0]),
            .clk                        (clk),
            .iwe                        (iwe));
      end
   endgenerate
endmodule


// Local Variables:
// verilog-library-directories:("." "sb_sim_rtl" )
// verilog-library-extensions:(".v" )
// End:
