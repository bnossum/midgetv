/* -----------------------------------------------------------------------------
 * Part of midgetv
 * 2019. Copyright B. Nossum.
 * For licence, see LICENCE
 * -----------------------------------------------------------------------------
 * EBR program memory is split into 2-bit wide memory, specified here.
 */
module m_ebr_w2
  # ( parameter [4095:0] prg0 = 4096'h0
      )
   (
    input [1:0]  B, //     Output from ALU
    input [10:0] Rai, //   Read adddress
    input [10:0] Wai, //   Write adddress
    input        clk, //   System clock
    input        we, //    Write enable
    output [1:0] DAT_O //  Registered output
    );

   /* verilator lint_off UNUSED */
   wire [13:0]   dum14;
   /* verilator lint_on UNUSED */

   SB_RAM40_4K 
     #(
       .INIT_F({prg0[4095],prg0[4093],prg0[4091],prg0[4089],prg0[4087],prg0[4085],prg0[4083],prg0[4081],
                prg0[4094],prg0[4092],prg0[4090],prg0[4088],prg0[4086],prg0[4084],prg0[4082],prg0[4080],
                prg0[4079],prg0[4077],prg0[4075],prg0[4073],prg0[4071],prg0[4069],prg0[4067],prg0[4065],
                prg0[4078],prg0[4076],prg0[4074],prg0[4072],prg0[4070],prg0[4068],prg0[4066],prg0[4064],
                prg0[4063],prg0[4061],prg0[4059],prg0[4057],prg0[4055],prg0[4053],prg0[4051],prg0[4049],
                prg0[4062],prg0[4060],prg0[4058],prg0[4056],prg0[4054],prg0[4052],prg0[4050],prg0[4048],
                prg0[4047],prg0[4045],prg0[4043],prg0[4041],prg0[4039],prg0[4037],prg0[4035],prg0[4033],
                prg0[4046],prg0[4044],prg0[4042],prg0[4040],prg0[4038],prg0[4036],prg0[4034],prg0[4032],
                prg0[4031],prg0[4029],prg0[4027],prg0[4025],prg0[4023],prg0[4021],prg0[4019],prg0[4017],
                prg0[4030],prg0[4028],prg0[4026],prg0[4024],prg0[4022],prg0[4020],prg0[4018],prg0[4016],
                prg0[4015],prg0[4013],prg0[4011],prg0[4009],prg0[4007],prg0[4005],prg0[4003],prg0[4001],
                prg0[4014],prg0[4012],prg0[4010],prg0[4008],prg0[4006],prg0[4004],prg0[4002],prg0[4000],
                prg0[3999],prg0[3997],prg0[3995],prg0[3993],prg0[3991],prg0[3989],prg0[3987],prg0[3985],
                prg0[3998],prg0[3996],prg0[3994],prg0[3992],prg0[3990],prg0[3988],prg0[3986],prg0[3984],
                prg0[3983],prg0[3981],prg0[3979],prg0[3977],prg0[3975],prg0[3973],prg0[3971],prg0[3969],
                prg0[3982],prg0[3980],prg0[3978],prg0[3976],prg0[3974],prg0[3972],prg0[3970],prg0[3968],
                prg0[3967],prg0[3965],prg0[3963],prg0[3961],prg0[3959],prg0[3957],prg0[3955],prg0[3953],
                prg0[3966],prg0[3964],prg0[3962],prg0[3960],prg0[3958],prg0[3956],prg0[3954],prg0[3952],
                prg0[3951],prg0[3949],prg0[3947],prg0[3945],prg0[3943],prg0[3941],prg0[3939],prg0[3937],
                prg0[3950],prg0[3948],prg0[3946],prg0[3944],prg0[3942],prg0[3940],prg0[3938],prg0[3936],
                prg0[3935],prg0[3933],prg0[3931],prg0[3929],prg0[3927],prg0[3925],prg0[3923],prg0[3921],
                prg0[3934],prg0[3932],prg0[3930],prg0[3928],prg0[3926],prg0[3924],prg0[3922],prg0[3920],
                prg0[3919],prg0[3917],prg0[3915],prg0[3913],prg0[3911],prg0[3909],prg0[3907],prg0[3905],
                prg0[3918],prg0[3916],prg0[3914],prg0[3912],prg0[3910],prg0[3908],prg0[3906],prg0[3904],
                prg0[3903],prg0[3901],prg0[3899],prg0[3897],prg0[3895],prg0[3893],prg0[3891],prg0[3889],
                prg0[3902],prg0[3900],prg0[3898],prg0[3896],prg0[3894],prg0[3892],prg0[3890],prg0[3888],
                prg0[3887],prg0[3885],prg0[3883],prg0[3881],prg0[3879],prg0[3877],prg0[3875],prg0[3873],
                prg0[3886],prg0[3884],prg0[3882],prg0[3880],prg0[3878],prg0[3876],prg0[3874],prg0[3872],
                prg0[3871],prg0[3869],prg0[3867],prg0[3865],prg0[3863],prg0[3861],prg0[3859],prg0[3857],
                prg0[3870],prg0[3868],prg0[3866],prg0[3864],prg0[3862],prg0[3860],prg0[3858],prg0[3856],
                prg0[3855],prg0[3853],prg0[3851],prg0[3849],prg0[3847],prg0[3845],prg0[3843],prg0[3841],
                prg0[3854],prg0[3852],prg0[3850],prg0[3848],prg0[3846],prg0[3844],prg0[3842],prg0[3840]}),
       .INIT_E({prg0[3839],prg0[3837],prg0[3835],prg0[3833],prg0[3831],prg0[3829],prg0[3827],prg0[3825],
                prg0[3838],prg0[3836],prg0[3834],prg0[3832],prg0[3830],prg0[3828],prg0[3826],prg0[3824],
                prg0[3823],prg0[3821],prg0[3819],prg0[3817],prg0[3815],prg0[3813],prg0[3811],prg0[3809],
                prg0[3822],prg0[3820],prg0[3818],prg0[3816],prg0[3814],prg0[3812],prg0[3810],prg0[3808],
                prg0[3807],prg0[3805],prg0[3803],prg0[3801],prg0[3799],prg0[3797],prg0[3795],prg0[3793],
                prg0[3806],prg0[3804],prg0[3802],prg0[3800],prg0[3798],prg0[3796],prg0[3794],prg0[3792],
                prg0[3791],prg0[3789],prg0[3787],prg0[3785],prg0[3783],prg0[3781],prg0[3779],prg0[3777],
                prg0[3790],prg0[3788],prg0[3786],prg0[3784],prg0[3782],prg0[3780],prg0[3778],prg0[3776],
                prg0[3775],prg0[3773],prg0[3771],prg0[3769],prg0[3767],prg0[3765],prg0[3763],prg0[3761],
                prg0[3774],prg0[3772],prg0[3770],prg0[3768],prg0[3766],prg0[3764],prg0[3762],prg0[3760],
                prg0[3759],prg0[3757],prg0[3755],prg0[3753],prg0[3751],prg0[3749],prg0[3747],prg0[3745],
                prg0[3758],prg0[3756],prg0[3754],prg0[3752],prg0[3750],prg0[3748],prg0[3746],prg0[3744],
                prg0[3743],prg0[3741],prg0[3739],prg0[3737],prg0[3735],prg0[3733],prg0[3731],prg0[3729],
                prg0[3742],prg0[3740],prg0[3738],prg0[3736],prg0[3734],prg0[3732],prg0[3730],prg0[3728],
                prg0[3727],prg0[3725],prg0[3723],prg0[3721],prg0[3719],prg0[3717],prg0[3715],prg0[3713],
                prg0[3726],prg0[3724],prg0[3722],prg0[3720],prg0[3718],prg0[3716],prg0[3714],prg0[3712],
                prg0[3711],prg0[3709],prg0[3707],prg0[3705],prg0[3703],prg0[3701],prg0[3699],prg0[3697],
                prg0[3710],prg0[3708],prg0[3706],prg0[3704],prg0[3702],prg0[3700],prg0[3698],prg0[3696],
                prg0[3695],prg0[3693],prg0[3691],prg0[3689],prg0[3687],prg0[3685],prg0[3683],prg0[3681],
                prg0[3694],prg0[3692],prg0[3690],prg0[3688],prg0[3686],prg0[3684],prg0[3682],prg0[3680],
                prg0[3679],prg0[3677],prg0[3675],prg0[3673],prg0[3671],prg0[3669],prg0[3667],prg0[3665],
                prg0[3678],prg0[3676],prg0[3674],prg0[3672],prg0[3670],prg0[3668],prg0[3666],prg0[3664],
                prg0[3663],prg0[3661],prg0[3659],prg0[3657],prg0[3655],prg0[3653],prg0[3651],prg0[3649],
                prg0[3662],prg0[3660],prg0[3658],prg0[3656],prg0[3654],prg0[3652],prg0[3650],prg0[3648],
                prg0[3647],prg0[3645],prg0[3643],prg0[3641],prg0[3639],prg0[3637],prg0[3635],prg0[3633],
                prg0[3646],prg0[3644],prg0[3642],prg0[3640],prg0[3638],prg0[3636],prg0[3634],prg0[3632],
                prg0[3631],prg0[3629],prg0[3627],prg0[3625],prg0[3623],prg0[3621],prg0[3619],prg0[3617],
                prg0[3630],prg0[3628],prg0[3626],prg0[3624],prg0[3622],prg0[3620],prg0[3618],prg0[3616],
                prg0[3615],prg0[3613],prg0[3611],prg0[3609],prg0[3607],prg0[3605],prg0[3603],prg0[3601],
                prg0[3614],prg0[3612],prg0[3610],prg0[3608],prg0[3606],prg0[3604],prg0[3602],prg0[3600],
                prg0[3599],prg0[3597],prg0[3595],prg0[3593],prg0[3591],prg0[3589],prg0[3587],prg0[3585],
                prg0[3598],prg0[3596],prg0[3594],prg0[3592],prg0[3590],prg0[3588],prg0[3586],prg0[3584]}),
       .INIT_D({prg0[3583],prg0[3581],prg0[3579],prg0[3577],prg0[3575],prg0[3573],prg0[3571],prg0[3569],
                prg0[3582],prg0[3580],prg0[3578],prg0[3576],prg0[3574],prg0[3572],prg0[3570],prg0[3568],
                prg0[3567],prg0[3565],prg0[3563],prg0[3561],prg0[3559],prg0[3557],prg0[3555],prg0[3553],
                prg0[3566],prg0[3564],prg0[3562],prg0[3560],prg0[3558],prg0[3556],prg0[3554],prg0[3552],
                prg0[3551],prg0[3549],prg0[3547],prg0[3545],prg0[3543],prg0[3541],prg0[3539],prg0[3537],
                prg0[3550],prg0[3548],prg0[3546],prg0[3544],prg0[3542],prg0[3540],prg0[3538],prg0[3536],
                prg0[3535],prg0[3533],prg0[3531],prg0[3529],prg0[3527],prg0[3525],prg0[3523],prg0[3521],
                prg0[3534],prg0[3532],prg0[3530],prg0[3528],prg0[3526],prg0[3524],prg0[3522],prg0[3520],
                prg0[3519],prg0[3517],prg0[3515],prg0[3513],prg0[3511],prg0[3509],prg0[3507],prg0[3505],
                prg0[3518],prg0[3516],prg0[3514],prg0[3512],prg0[3510],prg0[3508],prg0[3506],prg0[3504],
                prg0[3503],prg0[3501],prg0[3499],prg0[3497],prg0[3495],prg0[3493],prg0[3491],prg0[3489],
                prg0[3502],prg0[3500],prg0[3498],prg0[3496],prg0[3494],prg0[3492],prg0[3490],prg0[3488],
                prg0[3487],prg0[3485],prg0[3483],prg0[3481],prg0[3479],prg0[3477],prg0[3475],prg0[3473],
                prg0[3486],prg0[3484],prg0[3482],prg0[3480],prg0[3478],prg0[3476],prg0[3474],prg0[3472],
                prg0[3471],prg0[3469],prg0[3467],prg0[3465],prg0[3463],prg0[3461],prg0[3459],prg0[3457],
                prg0[3470],prg0[3468],prg0[3466],prg0[3464],prg0[3462],prg0[3460],prg0[3458],prg0[3456],
                prg0[3455],prg0[3453],prg0[3451],prg0[3449],prg0[3447],prg0[3445],prg0[3443],prg0[3441],
                prg0[3454],prg0[3452],prg0[3450],prg0[3448],prg0[3446],prg0[3444],prg0[3442],prg0[3440],
                prg0[3439],prg0[3437],prg0[3435],prg0[3433],prg0[3431],prg0[3429],prg0[3427],prg0[3425],
                prg0[3438],prg0[3436],prg0[3434],prg0[3432],prg0[3430],prg0[3428],prg0[3426],prg0[3424],
                prg0[3423],prg0[3421],prg0[3419],prg0[3417],prg0[3415],prg0[3413],prg0[3411],prg0[3409],
                prg0[3422],prg0[3420],prg0[3418],prg0[3416],prg0[3414],prg0[3412],prg0[3410],prg0[3408],
                prg0[3407],prg0[3405],prg0[3403],prg0[3401],prg0[3399],prg0[3397],prg0[3395],prg0[3393],
                prg0[3406],prg0[3404],prg0[3402],prg0[3400],prg0[3398],prg0[3396],prg0[3394],prg0[3392],
                prg0[3391],prg0[3389],prg0[3387],prg0[3385],prg0[3383],prg0[3381],prg0[3379],prg0[3377],
                prg0[3390],prg0[3388],prg0[3386],prg0[3384],prg0[3382],prg0[3380],prg0[3378],prg0[3376],
                prg0[3375],prg0[3373],prg0[3371],prg0[3369],prg0[3367],prg0[3365],prg0[3363],prg0[3361],
                prg0[3374],prg0[3372],prg0[3370],prg0[3368],prg0[3366],prg0[3364],prg0[3362],prg0[3360],
                prg0[3359],prg0[3357],prg0[3355],prg0[3353],prg0[3351],prg0[3349],prg0[3347],prg0[3345],
                prg0[3358],prg0[3356],prg0[3354],prg0[3352],prg0[3350],prg0[3348],prg0[3346],prg0[3344],
                prg0[3343],prg0[3341],prg0[3339],prg0[3337],prg0[3335],prg0[3333],prg0[3331],prg0[3329],
                prg0[3342],prg0[3340],prg0[3338],prg0[3336],prg0[3334],prg0[3332],prg0[3330],prg0[3328]}),
       .INIT_C({prg0[3327],prg0[3325],prg0[3323],prg0[3321],prg0[3319],prg0[3317],prg0[3315],prg0[3313],
                prg0[3326],prg0[3324],prg0[3322],prg0[3320],prg0[3318],prg0[3316],prg0[3314],prg0[3312],
                prg0[3311],prg0[3309],prg0[3307],prg0[3305],prg0[3303],prg0[3301],prg0[3299],prg0[3297],
                prg0[3310],prg0[3308],prg0[3306],prg0[3304],prg0[3302],prg0[3300],prg0[3298],prg0[3296],
                prg0[3295],prg0[3293],prg0[3291],prg0[3289],prg0[3287],prg0[3285],prg0[3283],prg0[3281],
                prg0[3294],prg0[3292],prg0[3290],prg0[3288],prg0[3286],prg0[3284],prg0[3282],prg0[3280],
                prg0[3279],prg0[3277],prg0[3275],prg0[3273],prg0[3271],prg0[3269],prg0[3267],prg0[3265],
                prg0[3278],prg0[3276],prg0[3274],prg0[3272],prg0[3270],prg0[3268],prg0[3266],prg0[3264],
                prg0[3263],prg0[3261],prg0[3259],prg0[3257],prg0[3255],prg0[3253],prg0[3251],prg0[3249],
                prg0[3262],prg0[3260],prg0[3258],prg0[3256],prg0[3254],prg0[3252],prg0[3250],prg0[3248],
                prg0[3247],prg0[3245],prg0[3243],prg0[3241],prg0[3239],prg0[3237],prg0[3235],prg0[3233],
                prg0[3246],prg0[3244],prg0[3242],prg0[3240],prg0[3238],prg0[3236],prg0[3234],prg0[3232],
                prg0[3231],prg0[3229],prg0[3227],prg0[3225],prg0[3223],prg0[3221],prg0[3219],prg0[3217],
                prg0[3230],prg0[3228],prg0[3226],prg0[3224],prg0[3222],prg0[3220],prg0[3218],prg0[3216],
                prg0[3215],prg0[3213],prg0[3211],prg0[3209],prg0[3207],prg0[3205],prg0[3203],prg0[3201],
                prg0[3214],prg0[3212],prg0[3210],prg0[3208],prg0[3206],prg0[3204],prg0[3202],prg0[3200],
                prg0[3199],prg0[3197],prg0[3195],prg0[3193],prg0[3191],prg0[3189],prg0[3187],prg0[3185],
                prg0[3198],prg0[3196],prg0[3194],prg0[3192],prg0[3190],prg0[3188],prg0[3186],prg0[3184],
                prg0[3183],prg0[3181],prg0[3179],prg0[3177],prg0[3175],prg0[3173],prg0[3171],prg0[3169],
                prg0[3182],prg0[3180],prg0[3178],prg0[3176],prg0[3174],prg0[3172],prg0[3170],prg0[3168],
                prg0[3167],prg0[3165],prg0[3163],prg0[3161],prg0[3159],prg0[3157],prg0[3155],prg0[3153],
                prg0[3166],prg0[3164],prg0[3162],prg0[3160],prg0[3158],prg0[3156],prg0[3154],prg0[3152],
                prg0[3151],prg0[3149],prg0[3147],prg0[3145],prg0[3143],prg0[3141],prg0[3139],prg0[3137],
                prg0[3150],prg0[3148],prg0[3146],prg0[3144],prg0[3142],prg0[3140],prg0[3138],prg0[3136],
                prg0[3135],prg0[3133],prg0[3131],prg0[3129],prg0[3127],prg0[3125],prg0[3123],prg0[3121],
                prg0[3134],prg0[3132],prg0[3130],prg0[3128],prg0[3126],prg0[3124],prg0[3122],prg0[3120],
                prg0[3119],prg0[3117],prg0[3115],prg0[3113],prg0[3111],prg0[3109],prg0[3107],prg0[3105],
                prg0[3118],prg0[3116],prg0[3114],prg0[3112],prg0[3110],prg0[3108],prg0[3106],prg0[3104],
                prg0[3103],prg0[3101],prg0[3099],prg0[3097],prg0[3095],prg0[3093],prg0[3091],prg0[3089],
                prg0[3102],prg0[3100],prg0[3098],prg0[3096],prg0[3094],prg0[3092],prg0[3090],prg0[3088],
                prg0[3087],prg0[3085],prg0[3083],prg0[3081],prg0[3079],prg0[3077],prg0[3075],prg0[3073],
                prg0[3086],prg0[3084],prg0[3082],prg0[3080],prg0[3078],prg0[3076],prg0[3074],prg0[3072]}),
       .INIT_B({prg0[3071],prg0[3069],prg0[3067],prg0[3065],prg0[3063],prg0[3061],prg0[3059],prg0[3057],
                prg0[3070],prg0[3068],prg0[3066],prg0[3064],prg0[3062],prg0[3060],prg0[3058],prg0[3056],
                prg0[3055],prg0[3053],prg0[3051],prg0[3049],prg0[3047],prg0[3045],prg0[3043],prg0[3041],
                prg0[3054],prg0[3052],prg0[3050],prg0[3048],prg0[3046],prg0[3044],prg0[3042],prg0[3040],
                prg0[3039],prg0[3037],prg0[3035],prg0[3033],prg0[3031],prg0[3029],prg0[3027],prg0[3025],
                prg0[3038],prg0[3036],prg0[3034],prg0[3032],prg0[3030],prg0[3028],prg0[3026],prg0[3024],
                prg0[3023],prg0[3021],prg0[3019],prg0[3017],prg0[3015],prg0[3013],prg0[3011],prg0[3009],
                prg0[3022],prg0[3020],prg0[3018],prg0[3016],prg0[3014],prg0[3012],prg0[3010],prg0[3008],
                prg0[3007],prg0[3005],prg0[3003],prg0[3001],prg0[2999],prg0[2997],prg0[2995],prg0[2993],
                prg0[3006],prg0[3004],prg0[3002],prg0[3000],prg0[2998],prg0[2996],prg0[2994],prg0[2992],
                prg0[2991],prg0[2989],prg0[2987],prg0[2985],prg0[2983],prg0[2981],prg0[2979],prg0[2977],
                prg0[2990],prg0[2988],prg0[2986],prg0[2984],prg0[2982],prg0[2980],prg0[2978],prg0[2976],
                prg0[2975],prg0[2973],prg0[2971],prg0[2969],prg0[2967],prg0[2965],prg0[2963],prg0[2961],
                prg0[2974],prg0[2972],prg0[2970],prg0[2968],prg0[2966],prg0[2964],prg0[2962],prg0[2960],
                prg0[2959],prg0[2957],prg0[2955],prg0[2953],prg0[2951],prg0[2949],prg0[2947],prg0[2945],
                prg0[2958],prg0[2956],prg0[2954],prg0[2952],prg0[2950],prg0[2948],prg0[2946],prg0[2944],
                prg0[2943],prg0[2941],prg0[2939],prg0[2937],prg0[2935],prg0[2933],prg0[2931],prg0[2929],
                prg0[2942],prg0[2940],prg0[2938],prg0[2936],prg0[2934],prg0[2932],prg0[2930],prg0[2928],
                prg0[2927],prg0[2925],prg0[2923],prg0[2921],prg0[2919],prg0[2917],prg0[2915],prg0[2913],
                prg0[2926],prg0[2924],prg0[2922],prg0[2920],prg0[2918],prg0[2916],prg0[2914],prg0[2912],
                prg0[2911],prg0[2909],prg0[2907],prg0[2905],prg0[2903],prg0[2901],prg0[2899],prg0[2897],
                prg0[2910],prg0[2908],prg0[2906],prg0[2904],prg0[2902],prg0[2900],prg0[2898],prg0[2896],
                prg0[2895],prg0[2893],prg0[2891],prg0[2889],prg0[2887],prg0[2885],prg0[2883],prg0[2881],
                prg0[2894],prg0[2892],prg0[2890],prg0[2888],prg0[2886],prg0[2884],prg0[2882],prg0[2880],
                prg0[2879],prg0[2877],prg0[2875],prg0[2873],prg0[2871],prg0[2869],prg0[2867],prg0[2865],
                prg0[2878],prg0[2876],prg0[2874],prg0[2872],prg0[2870],prg0[2868],prg0[2866],prg0[2864],
                prg0[2863],prg0[2861],prg0[2859],prg0[2857],prg0[2855],prg0[2853],prg0[2851],prg0[2849],
                prg0[2862],prg0[2860],prg0[2858],prg0[2856],prg0[2854],prg0[2852],prg0[2850],prg0[2848],
                prg0[2847],prg0[2845],prg0[2843],prg0[2841],prg0[2839],prg0[2837],prg0[2835],prg0[2833],
                prg0[2846],prg0[2844],prg0[2842],prg0[2840],prg0[2838],prg0[2836],prg0[2834],prg0[2832],
                prg0[2831],prg0[2829],prg0[2827],prg0[2825],prg0[2823],prg0[2821],prg0[2819],prg0[2817],
                prg0[2830],prg0[2828],prg0[2826],prg0[2824],prg0[2822],prg0[2820],prg0[2818],prg0[2816]}),
       .INIT_A({prg0[2815],prg0[2813],prg0[2811],prg0[2809],prg0[2807],prg0[2805],prg0[2803],prg0[2801],
                prg0[2814],prg0[2812],prg0[2810],prg0[2808],prg0[2806],prg0[2804],prg0[2802],prg0[2800],
                prg0[2799],prg0[2797],prg0[2795],prg0[2793],prg0[2791],prg0[2789],prg0[2787],prg0[2785],
                prg0[2798],prg0[2796],prg0[2794],prg0[2792],prg0[2790],prg0[2788],prg0[2786],prg0[2784],
                prg0[2783],prg0[2781],prg0[2779],prg0[2777],prg0[2775],prg0[2773],prg0[2771],prg0[2769],
                prg0[2782],prg0[2780],prg0[2778],prg0[2776],prg0[2774],prg0[2772],prg0[2770],prg0[2768],
                prg0[2767],prg0[2765],prg0[2763],prg0[2761],prg0[2759],prg0[2757],prg0[2755],prg0[2753],
                prg0[2766],prg0[2764],prg0[2762],prg0[2760],prg0[2758],prg0[2756],prg0[2754],prg0[2752],
                prg0[2751],prg0[2749],prg0[2747],prg0[2745],prg0[2743],prg0[2741],prg0[2739],prg0[2737],
                prg0[2750],prg0[2748],prg0[2746],prg0[2744],prg0[2742],prg0[2740],prg0[2738],prg0[2736],
                prg0[2735],prg0[2733],prg0[2731],prg0[2729],prg0[2727],prg0[2725],prg0[2723],prg0[2721],
                prg0[2734],prg0[2732],prg0[2730],prg0[2728],prg0[2726],prg0[2724],prg0[2722],prg0[2720],
                prg0[2719],prg0[2717],prg0[2715],prg0[2713],prg0[2711],prg0[2709],prg0[2707],prg0[2705],
                prg0[2718],prg0[2716],prg0[2714],prg0[2712],prg0[2710],prg0[2708],prg0[2706],prg0[2704],
                prg0[2703],prg0[2701],prg0[2699],prg0[2697],prg0[2695],prg0[2693],prg0[2691],prg0[2689],
                prg0[2702],prg0[2700],prg0[2698],prg0[2696],prg0[2694],prg0[2692],prg0[2690],prg0[2688],
                prg0[2687],prg0[2685],prg0[2683],prg0[2681],prg0[2679],prg0[2677],prg0[2675],prg0[2673],
                prg0[2686],prg0[2684],prg0[2682],prg0[2680],prg0[2678],prg0[2676],prg0[2674],prg0[2672],
                prg0[2671],prg0[2669],prg0[2667],prg0[2665],prg0[2663],prg0[2661],prg0[2659],prg0[2657],
                prg0[2670],prg0[2668],prg0[2666],prg0[2664],prg0[2662],prg0[2660],prg0[2658],prg0[2656],
                prg0[2655],prg0[2653],prg0[2651],prg0[2649],prg0[2647],prg0[2645],prg0[2643],prg0[2641],
                prg0[2654],prg0[2652],prg0[2650],prg0[2648],prg0[2646],prg0[2644],prg0[2642],prg0[2640],
                prg0[2639],prg0[2637],prg0[2635],prg0[2633],prg0[2631],prg0[2629],prg0[2627],prg0[2625],
                prg0[2638],prg0[2636],prg0[2634],prg0[2632],prg0[2630],prg0[2628],prg0[2626],prg0[2624],
                prg0[2623],prg0[2621],prg0[2619],prg0[2617],prg0[2615],prg0[2613],prg0[2611],prg0[2609],
                prg0[2622],prg0[2620],prg0[2618],prg0[2616],prg0[2614],prg0[2612],prg0[2610],prg0[2608],
                prg0[2607],prg0[2605],prg0[2603],prg0[2601],prg0[2599],prg0[2597],prg0[2595],prg0[2593],
                prg0[2606],prg0[2604],prg0[2602],prg0[2600],prg0[2598],prg0[2596],prg0[2594],prg0[2592],
                prg0[2591],prg0[2589],prg0[2587],prg0[2585],prg0[2583],prg0[2581],prg0[2579],prg0[2577],
                prg0[2590],prg0[2588],prg0[2586],prg0[2584],prg0[2582],prg0[2580],prg0[2578],prg0[2576],
                prg0[2575],prg0[2573],prg0[2571],prg0[2569],prg0[2567],prg0[2565],prg0[2563],prg0[2561],
                prg0[2574],prg0[2572],prg0[2570],prg0[2568],prg0[2566],prg0[2564],prg0[2562],prg0[2560]}),
       .INIT_9({prg0[2559],prg0[2557],prg0[2555],prg0[2553],prg0[2551],prg0[2549],prg0[2547],prg0[2545],
                prg0[2558],prg0[2556],prg0[2554],prg0[2552],prg0[2550],prg0[2548],prg0[2546],prg0[2544],
                prg0[2543],prg0[2541],prg0[2539],prg0[2537],prg0[2535],prg0[2533],prg0[2531],prg0[2529],
                prg0[2542],prg0[2540],prg0[2538],prg0[2536],prg0[2534],prg0[2532],prg0[2530],prg0[2528],
                prg0[2527],prg0[2525],prg0[2523],prg0[2521],prg0[2519],prg0[2517],prg0[2515],prg0[2513],
                prg0[2526],prg0[2524],prg0[2522],prg0[2520],prg0[2518],prg0[2516],prg0[2514],prg0[2512],
                prg0[2511],prg0[2509],prg0[2507],prg0[2505],prg0[2503],prg0[2501],prg0[2499],prg0[2497],
                prg0[2510],prg0[2508],prg0[2506],prg0[2504],prg0[2502],prg0[2500],prg0[2498],prg0[2496],
                prg0[2495],prg0[2493],prg0[2491],prg0[2489],prg0[2487],prg0[2485],prg0[2483],prg0[2481],
                prg0[2494],prg0[2492],prg0[2490],prg0[2488],prg0[2486],prg0[2484],prg0[2482],prg0[2480],
                prg0[2479],prg0[2477],prg0[2475],prg0[2473],prg0[2471],prg0[2469],prg0[2467],prg0[2465],
                prg0[2478],prg0[2476],prg0[2474],prg0[2472],prg0[2470],prg0[2468],prg0[2466],prg0[2464],
                prg0[2463],prg0[2461],prg0[2459],prg0[2457],prg0[2455],prg0[2453],prg0[2451],prg0[2449],
                prg0[2462],prg0[2460],prg0[2458],prg0[2456],prg0[2454],prg0[2452],prg0[2450],prg0[2448],
                prg0[2447],prg0[2445],prg0[2443],prg0[2441],prg0[2439],prg0[2437],prg0[2435],prg0[2433],
                prg0[2446],prg0[2444],prg0[2442],prg0[2440],prg0[2438],prg0[2436],prg0[2434],prg0[2432],
                prg0[2431],prg0[2429],prg0[2427],prg0[2425],prg0[2423],prg0[2421],prg0[2419],prg0[2417],
                prg0[2430],prg0[2428],prg0[2426],prg0[2424],prg0[2422],prg0[2420],prg0[2418],prg0[2416],
                prg0[2415],prg0[2413],prg0[2411],prg0[2409],prg0[2407],prg0[2405],prg0[2403],prg0[2401],
                prg0[2414],prg0[2412],prg0[2410],prg0[2408],prg0[2406],prg0[2404],prg0[2402],prg0[2400],
                prg0[2399],prg0[2397],prg0[2395],prg0[2393],prg0[2391],prg0[2389],prg0[2387],prg0[2385],
                prg0[2398],prg0[2396],prg0[2394],prg0[2392],prg0[2390],prg0[2388],prg0[2386],prg0[2384],
                prg0[2383],prg0[2381],prg0[2379],prg0[2377],prg0[2375],prg0[2373],prg0[2371],prg0[2369],
                prg0[2382],prg0[2380],prg0[2378],prg0[2376],prg0[2374],prg0[2372],prg0[2370],prg0[2368],
                prg0[2367],prg0[2365],prg0[2363],prg0[2361],prg0[2359],prg0[2357],prg0[2355],prg0[2353],
                prg0[2366],prg0[2364],prg0[2362],prg0[2360],prg0[2358],prg0[2356],prg0[2354],prg0[2352],
                prg0[2351],prg0[2349],prg0[2347],prg0[2345],prg0[2343],prg0[2341],prg0[2339],prg0[2337],
                prg0[2350],prg0[2348],prg0[2346],prg0[2344],prg0[2342],prg0[2340],prg0[2338],prg0[2336],
                prg0[2335],prg0[2333],prg0[2331],prg0[2329],prg0[2327],prg0[2325],prg0[2323],prg0[2321],
                prg0[2334],prg0[2332],prg0[2330],prg0[2328],prg0[2326],prg0[2324],prg0[2322],prg0[2320],
                prg0[2319],prg0[2317],prg0[2315],prg0[2313],prg0[2311],prg0[2309],prg0[2307],prg0[2305],
                prg0[2318],prg0[2316],prg0[2314],prg0[2312],prg0[2310],prg0[2308],prg0[2306],prg0[2304]}),
       .INIT_8({prg0[2303],prg0[2301],prg0[2299],prg0[2297],prg0[2295],prg0[2293],prg0[2291],prg0[2289],
                prg0[2302],prg0[2300],prg0[2298],prg0[2296],prg0[2294],prg0[2292],prg0[2290],prg0[2288],
                prg0[2287],prg0[2285],prg0[2283],prg0[2281],prg0[2279],prg0[2277],prg0[2275],prg0[2273],
                prg0[2286],prg0[2284],prg0[2282],prg0[2280],prg0[2278],prg0[2276],prg0[2274],prg0[2272],
                prg0[2271],prg0[2269],prg0[2267],prg0[2265],prg0[2263],prg0[2261],prg0[2259],prg0[2257],
                prg0[2270],prg0[2268],prg0[2266],prg0[2264],prg0[2262],prg0[2260],prg0[2258],prg0[2256],
                prg0[2255],prg0[2253],prg0[2251],prg0[2249],prg0[2247],prg0[2245],prg0[2243],prg0[2241],
                prg0[2254],prg0[2252],prg0[2250],prg0[2248],prg0[2246],prg0[2244],prg0[2242],prg0[2240],
                prg0[2239],prg0[2237],prg0[2235],prg0[2233],prg0[2231],prg0[2229],prg0[2227],prg0[2225],
                prg0[2238],prg0[2236],prg0[2234],prg0[2232],prg0[2230],prg0[2228],prg0[2226],prg0[2224],
                prg0[2223],prg0[2221],prg0[2219],prg0[2217],prg0[2215],prg0[2213],prg0[2211],prg0[2209],
                prg0[2222],prg0[2220],prg0[2218],prg0[2216],prg0[2214],prg0[2212],prg0[2210],prg0[2208],
                prg0[2207],prg0[2205],prg0[2203],prg0[2201],prg0[2199],prg0[2197],prg0[2195],prg0[2193],
                prg0[2206],prg0[2204],prg0[2202],prg0[2200],prg0[2198],prg0[2196],prg0[2194],prg0[2192],
                prg0[2191],prg0[2189],prg0[2187],prg0[2185],prg0[2183],prg0[2181],prg0[2179],prg0[2177],
                prg0[2190],prg0[2188],prg0[2186],prg0[2184],prg0[2182],prg0[2180],prg0[2178],prg0[2176],
                prg0[2175],prg0[2173],prg0[2171],prg0[2169],prg0[2167],prg0[2165],prg0[2163],prg0[2161],
                prg0[2174],prg0[2172],prg0[2170],prg0[2168],prg0[2166],prg0[2164],prg0[2162],prg0[2160],
                prg0[2159],prg0[2157],prg0[2155],prg0[2153],prg0[2151],prg0[2149],prg0[2147],prg0[2145],
                prg0[2158],prg0[2156],prg0[2154],prg0[2152],prg0[2150],prg0[2148],prg0[2146],prg0[2144],
                prg0[2143],prg0[2141],prg0[2139],prg0[2137],prg0[2135],prg0[2133],prg0[2131],prg0[2129],
                prg0[2142],prg0[2140],prg0[2138],prg0[2136],prg0[2134],prg0[2132],prg0[2130],prg0[2128],
                prg0[2127],prg0[2125],prg0[2123],prg0[2121],prg0[2119],prg0[2117],prg0[2115],prg0[2113],
                prg0[2126],prg0[2124],prg0[2122],prg0[2120],prg0[2118],prg0[2116],prg0[2114],prg0[2112],
                prg0[2111],prg0[2109],prg0[2107],prg0[2105],prg0[2103],prg0[2101],prg0[2099],prg0[2097],
                prg0[2110],prg0[2108],prg0[2106],prg0[2104],prg0[2102],prg0[2100],prg0[2098],prg0[2096],
                prg0[2095],prg0[2093],prg0[2091],prg0[2089],prg0[2087],prg0[2085],prg0[2083],prg0[2081],
                prg0[2094],prg0[2092],prg0[2090],prg0[2088],prg0[2086],prg0[2084],prg0[2082],prg0[2080],
                prg0[2079],prg0[2077],prg0[2075],prg0[2073],prg0[2071],prg0[2069],prg0[2067],prg0[2065],
                prg0[2078],prg0[2076],prg0[2074],prg0[2072],prg0[2070],prg0[2068],prg0[2066],prg0[2064],
                prg0[2063],prg0[2061],prg0[2059],prg0[2057],prg0[2055],prg0[2053],prg0[2051],prg0[2049],
                prg0[2062],prg0[2060],prg0[2058],prg0[2056],prg0[2054],prg0[2052],prg0[2050],prg0[2048]}),
       .INIT_7({prg0[2047],prg0[2045],prg0[2043],prg0[2041],prg0[2039],prg0[2037],prg0[2035],prg0[2033],
                prg0[2046],prg0[2044],prg0[2042],prg0[2040],prg0[2038],prg0[2036],prg0[2034],prg0[2032],
                prg0[2031],prg0[2029],prg0[2027],prg0[2025],prg0[2023],prg0[2021],prg0[2019],prg0[2017],
                prg0[2030],prg0[2028],prg0[2026],prg0[2024],prg0[2022],prg0[2020],prg0[2018],prg0[2016],
                prg0[2015],prg0[2013],prg0[2011],prg0[2009],prg0[2007],prg0[2005],prg0[2003],prg0[2001],
                prg0[2014],prg0[2012],prg0[2010],prg0[2008],prg0[2006],prg0[2004],prg0[2002],prg0[2000],
                prg0[1999],prg0[1997],prg0[1995],prg0[1993],prg0[1991],prg0[1989],prg0[1987],prg0[1985],
                prg0[1998],prg0[1996],prg0[1994],prg0[1992],prg0[1990],prg0[1988],prg0[1986],prg0[1984],
                prg0[1983],prg0[1981],prg0[1979],prg0[1977],prg0[1975],prg0[1973],prg0[1971],prg0[1969],
                prg0[1982],prg0[1980],prg0[1978],prg0[1976],prg0[1974],prg0[1972],prg0[1970],prg0[1968],
                prg0[1967],prg0[1965],prg0[1963],prg0[1961],prg0[1959],prg0[1957],prg0[1955],prg0[1953],
                prg0[1966],prg0[1964],prg0[1962],prg0[1960],prg0[1958],prg0[1956],prg0[1954],prg0[1952],
                prg0[1951],prg0[1949],prg0[1947],prg0[1945],prg0[1943],prg0[1941],prg0[1939],prg0[1937],
                prg0[1950],prg0[1948],prg0[1946],prg0[1944],prg0[1942],prg0[1940],prg0[1938],prg0[1936],
                prg0[1935],prg0[1933],prg0[1931],prg0[1929],prg0[1927],prg0[1925],prg0[1923],prg0[1921],
                prg0[1934],prg0[1932],prg0[1930],prg0[1928],prg0[1926],prg0[1924],prg0[1922],prg0[1920],
                prg0[1919],prg0[1917],prg0[1915],prg0[1913],prg0[1911],prg0[1909],prg0[1907],prg0[1905],
                prg0[1918],prg0[1916],prg0[1914],prg0[1912],prg0[1910],prg0[1908],prg0[1906],prg0[1904],
                prg0[1903],prg0[1901],prg0[1899],prg0[1897],prg0[1895],prg0[1893],prg0[1891],prg0[1889],
                prg0[1902],prg0[1900],prg0[1898],prg0[1896],prg0[1894],prg0[1892],prg0[1890],prg0[1888],
                prg0[1887],prg0[1885],prg0[1883],prg0[1881],prg0[1879],prg0[1877],prg0[1875],prg0[1873],
                prg0[1886],prg0[1884],prg0[1882],prg0[1880],prg0[1878],prg0[1876],prg0[1874],prg0[1872],
                prg0[1871],prg0[1869],prg0[1867],prg0[1865],prg0[1863],prg0[1861],prg0[1859],prg0[1857],
                prg0[1870],prg0[1868],prg0[1866],prg0[1864],prg0[1862],prg0[1860],prg0[1858],prg0[1856],
                prg0[1855],prg0[1853],prg0[1851],prg0[1849],prg0[1847],prg0[1845],prg0[1843],prg0[1841],
                prg0[1854],prg0[1852],prg0[1850],prg0[1848],prg0[1846],prg0[1844],prg0[1842],prg0[1840],
                prg0[1839],prg0[1837],prg0[1835],prg0[1833],prg0[1831],prg0[1829],prg0[1827],prg0[1825],
                prg0[1838],prg0[1836],prg0[1834],prg0[1832],prg0[1830],prg0[1828],prg0[1826],prg0[1824],
                prg0[1823],prg0[1821],prg0[1819],prg0[1817],prg0[1815],prg0[1813],prg0[1811],prg0[1809],
                prg0[1822],prg0[1820],prg0[1818],prg0[1816],prg0[1814],prg0[1812],prg0[1810],prg0[1808],
                prg0[1807],prg0[1805],prg0[1803],prg0[1801],prg0[1799],prg0[1797],prg0[1795],prg0[1793],
                prg0[1806],prg0[1804],prg0[1802],prg0[1800],prg0[1798],prg0[1796],prg0[1794],prg0[1792]}),
       .INIT_6({prg0[1791],prg0[1789],prg0[1787],prg0[1785],prg0[1783],prg0[1781],prg0[1779],prg0[1777],
                prg0[1790],prg0[1788],prg0[1786],prg0[1784],prg0[1782],prg0[1780],prg0[1778],prg0[1776],
                prg0[1775],prg0[1773],prg0[1771],prg0[1769],prg0[1767],prg0[1765],prg0[1763],prg0[1761],
                prg0[1774],prg0[1772],prg0[1770],prg0[1768],prg0[1766],prg0[1764],prg0[1762],prg0[1760],
                prg0[1759],prg0[1757],prg0[1755],prg0[1753],prg0[1751],prg0[1749],prg0[1747],prg0[1745],
                prg0[1758],prg0[1756],prg0[1754],prg0[1752],prg0[1750],prg0[1748],prg0[1746],prg0[1744],
                prg0[1743],prg0[1741],prg0[1739],prg0[1737],prg0[1735],prg0[1733],prg0[1731],prg0[1729],
                prg0[1742],prg0[1740],prg0[1738],prg0[1736],prg0[1734],prg0[1732],prg0[1730],prg0[1728],
                prg0[1727],prg0[1725],prg0[1723],prg0[1721],prg0[1719],prg0[1717],prg0[1715],prg0[1713],
                prg0[1726],prg0[1724],prg0[1722],prg0[1720],prg0[1718],prg0[1716],prg0[1714],prg0[1712],
                prg0[1711],prg0[1709],prg0[1707],prg0[1705],prg0[1703],prg0[1701],prg0[1699],prg0[1697],
                prg0[1710],prg0[1708],prg0[1706],prg0[1704],prg0[1702],prg0[1700],prg0[1698],prg0[1696],
                prg0[1695],prg0[1693],prg0[1691],prg0[1689],prg0[1687],prg0[1685],prg0[1683],prg0[1681],
                prg0[1694],prg0[1692],prg0[1690],prg0[1688],prg0[1686],prg0[1684],prg0[1682],prg0[1680],
                prg0[1679],prg0[1677],prg0[1675],prg0[1673],prg0[1671],prg0[1669],prg0[1667],prg0[1665],
                prg0[1678],prg0[1676],prg0[1674],prg0[1672],prg0[1670],prg0[1668],prg0[1666],prg0[1664],
                prg0[1663],prg0[1661],prg0[1659],prg0[1657],prg0[1655],prg0[1653],prg0[1651],prg0[1649],
                prg0[1662],prg0[1660],prg0[1658],prg0[1656],prg0[1654],prg0[1652],prg0[1650],prg0[1648],
                prg0[1647],prg0[1645],prg0[1643],prg0[1641],prg0[1639],prg0[1637],prg0[1635],prg0[1633],
                prg0[1646],prg0[1644],prg0[1642],prg0[1640],prg0[1638],prg0[1636],prg0[1634],prg0[1632],
                prg0[1631],prg0[1629],prg0[1627],prg0[1625],prg0[1623],prg0[1621],prg0[1619],prg0[1617],
                prg0[1630],prg0[1628],prg0[1626],prg0[1624],prg0[1622],prg0[1620],prg0[1618],prg0[1616],
                prg0[1615],prg0[1613],prg0[1611],prg0[1609],prg0[1607],prg0[1605],prg0[1603],prg0[1601],
                prg0[1614],prg0[1612],prg0[1610],prg0[1608],prg0[1606],prg0[1604],prg0[1602],prg0[1600],
                prg0[1599],prg0[1597],prg0[1595],prg0[1593],prg0[1591],prg0[1589],prg0[1587],prg0[1585],
                prg0[1598],prg0[1596],prg0[1594],prg0[1592],prg0[1590],prg0[1588],prg0[1586],prg0[1584],
                prg0[1583],prg0[1581],prg0[1579],prg0[1577],prg0[1575],prg0[1573],prg0[1571],prg0[1569],
                prg0[1582],prg0[1580],prg0[1578],prg0[1576],prg0[1574],prg0[1572],prg0[1570],prg0[1568],
                prg0[1567],prg0[1565],prg0[1563],prg0[1561],prg0[1559],prg0[1557],prg0[1555],prg0[1553],
                prg0[1566],prg0[1564],prg0[1562],prg0[1560],prg0[1558],prg0[1556],prg0[1554],prg0[1552],
                prg0[1551],prg0[1549],prg0[1547],prg0[1545],prg0[1543],prg0[1541],prg0[1539],prg0[1537],
                prg0[1550],prg0[1548],prg0[1546],prg0[1544],prg0[1542],prg0[1540],prg0[1538],prg0[1536]}),
       .INIT_5({prg0[1535],prg0[1533],prg0[1531],prg0[1529],prg0[1527],prg0[1525],prg0[1523],prg0[1521],
                prg0[1534],prg0[1532],prg0[1530],prg0[1528],prg0[1526],prg0[1524],prg0[1522],prg0[1520],
                prg0[1519],prg0[1517],prg0[1515],prg0[1513],prg0[1511],prg0[1509],prg0[1507],prg0[1505],
                prg0[1518],prg0[1516],prg0[1514],prg0[1512],prg0[1510],prg0[1508],prg0[1506],prg0[1504],
                prg0[1503],prg0[1501],prg0[1499],prg0[1497],prg0[1495],prg0[1493],prg0[1491],prg0[1489],
                prg0[1502],prg0[1500],prg0[1498],prg0[1496],prg0[1494],prg0[1492],prg0[1490],prg0[1488],
                prg0[1487],prg0[1485],prg0[1483],prg0[1481],prg0[1479],prg0[1477],prg0[1475],prg0[1473],
                prg0[1486],prg0[1484],prg0[1482],prg0[1480],prg0[1478],prg0[1476],prg0[1474],prg0[1472],
                prg0[1471],prg0[1469],prg0[1467],prg0[1465],prg0[1463],prg0[1461],prg0[1459],prg0[1457],
                prg0[1470],prg0[1468],prg0[1466],prg0[1464],prg0[1462],prg0[1460],prg0[1458],prg0[1456],
                prg0[1455],prg0[1453],prg0[1451],prg0[1449],prg0[1447],prg0[1445],prg0[1443],prg0[1441],
                prg0[1454],prg0[1452],prg0[1450],prg0[1448],prg0[1446],prg0[1444],prg0[1442],prg0[1440],
                prg0[1439],prg0[1437],prg0[1435],prg0[1433],prg0[1431],prg0[1429],prg0[1427],prg0[1425],
                prg0[1438],prg0[1436],prg0[1434],prg0[1432],prg0[1430],prg0[1428],prg0[1426],prg0[1424],
                prg0[1423],prg0[1421],prg0[1419],prg0[1417],prg0[1415],prg0[1413],prg0[1411],prg0[1409],
                prg0[1422],prg0[1420],prg0[1418],prg0[1416],prg0[1414],prg0[1412],prg0[1410],prg0[1408],
                prg0[1407],prg0[1405],prg0[1403],prg0[1401],prg0[1399],prg0[1397],prg0[1395],prg0[1393],
                prg0[1406],prg0[1404],prg0[1402],prg0[1400],prg0[1398],prg0[1396],prg0[1394],prg0[1392],
                prg0[1391],prg0[1389],prg0[1387],prg0[1385],prg0[1383],prg0[1381],prg0[1379],prg0[1377],
                prg0[1390],prg0[1388],prg0[1386],prg0[1384],prg0[1382],prg0[1380],prg0[1378],prg0[1376],
                prg0[1375],prg0[1373],prg0[1371],prg0[1369],prg0[1367],prg0[1365],prg0[1363],prg0[1361],
                prg0[1374],prg0[1372],prg0[1370],prg0[1368],prg0[1366],prg0[1364],prg0[1362],prg0[1360],
                prg0[1359],prg0[1357],prg0[1355],prg0[1353],prg0[1351],prg0[1349],prg0[1347],prg0[1345],
                prg0[1358],prg0[1356],prg0[1354],prg0[1352],prg0[1350],prg0[1348],prg0[1346],prg0[1344],
                prg0[1343],prg0[1341],prg0[1339],prg0[1337],prg0[1335],prg0[1333],prg0[1331],prg0[1329],
                prg0[1342],prg0[1340],prg0[1338],prg0[1336],prg0[1334],prg0[1332],prg0[1330],prg0[1328],
                prg0[1327],prg0[1325],prg0[1323],prg0[1321],prg0[1319],prg0[1317],prg0[1315],prg0[1313],
                prg0[1326],prg0[1324],prg0[1322],prg0[1320],prg0[1318],prg0[1316],prg0[1314],prg0[1312],
                prg0[1311],prg0[1309],prg0[1307],prg0[1305],prg0[1303],prg0[1301],prg0[1299],prg0[1297],
                prg0[1310],prg0[1308],prg0[1306],prg0[1304],prg0[1302],prg0[1300],prg0[1298],prg0[1296],
                prg0[1295],prg0[1293],prg0[1291],prg0[1289],prg0[1287],prg0[1285],prg0[1283],prg0[1281],
                prg0[1294],prg0[1292],prg0[1290],prg0[1288],prg0[1286],prg0[1284],prg0[1282],prg0[1280]}),
       .INIT_4({prg0[1279],prg0[1277],prg0[1275],prg0[1273],prg0[1271],prg0[1269],prg0[1267],prg0[1265],
                prg0[1278],prg0[1276],prg0[1274],prg0[1272],prg0[1270],prg0[1268],prg0[1266],prg0[1264],
                prg0[1263],prg0[1261],prg0[1259],prg0[1257],prg0[1255],prg0[1253],prg0[1251],prg0[1249],
                prg0[1262],prg0[1260],prg0[1258],prg0[1256],prg0[1254],prg0[1252],prg0[1250],prg0[1248],
                prg0[1247],prg0[1245],prg0[1243],prg0[1241],prg0[1239],prg0[1237],prg0[1235],prg0[1233],
                prg0[1246],prg0[1244],prg0[1242],prg0[1240],prg0[1238],prg0[1236],prg0[1234],prg0[1232],
                prg0[1231],prg0[1229],prg0[1227],prg0[1225],prg0[1223],prg0[1221],prg0[1219],prg0[1217],
                prg0[1230],prg0[1228],prg0[1226],prg0[1224],prg0[1222],prg0[1220],prg0[1218],prg0[1216],
                prg0[1215],prg0[1213],prg0[1211],prg0[1209],prg0[1207],prg0[1205],prg0[1203],prg0[1201],
                prg0[1214],prg0[1212],prg0[1210],prg0[1208],prg0[1206],prg0[1204],prg0[1202],prg0[1200],
                prg0[1199],prg0[1197],prg0[1195],prg0[1193],prg0[1191],prg0[1189],prg0[1187],prg0[1185],
                prg0[1198],prg0[1196],prg0[1194],prg0[1192],prg0[1190],prg0[1188],prg0[1186],prg0[1184],
                prg0[1183],prg0[1181],prg0[1179],prg0[1177],prg0[1175],prg0[1173],prg0[1171],prg0[1169],
                prg0[1182],prg0[1180],prg0[1178],prg0[1176],prg0[1174],prg0[1172],prg0[1170],prg0[1168],
                prg0[1167],prg0[1165],prg0[1163],prg0[1161],prg0[1159],prg0[1157],prg0[1155],prg0[1153],
                prg0[1166],prg0[1164],prg0[1162],prg0[1160],prg0[1158],prg0[1156],prg0[1154],prg0[1152],
                prg0[1151],prg0[1149],prg0[1147],prg0[1145],prg0[1143],prg0[1141],prg0[1139],prg0[1137],
                prg0[1150],prg0[1148],prg0[1146],prg0[1144],prg0[1142],prg0[1140],prg0[1138],prg0[1136],
                prg0[1135],prg0[1133],prg0[1131],prg0[1129],prg0[1127],prg0[1125],prg0[1123],prg0[1121],
                prg0[1134],prg0[1132],prg0[1130],prg0[1128],prg0[1126],prg0[1124],prg0[1122],prg0[1120],
                prg0[1119],prg0[1117],prg0[1115],prg0[1113],prg0[1111],prg0[1109],prg0[1107],prg0[1105],
                prg0[1118],prg0[1116],prg0[1114],prg0[1112],prg0[1110],prg0[1108],prg0[1106],prg0[1104],
                prg0[1103],prg0[1101],prg0[1099],prg0[1097],prg0[1095],prg0[1093],prg0[1091],prg0[1089],
                prg0[1102],prg0[1100],prg0[1098],prg0[1096],prg0[1094],prg0[1092],prg0[1090],prg0[1088],
                prg0[1087],prg0[1085],prg0[1083],prg0[1081],prg0[1079],prg0[1077],prg0[1075],prg0[1073],
                prg0[1086],prg0[1084],prg0[1082],prg0[1080],prg0[1078],prg0[1076],prg0[1074],prg0[1072],
                prg0[1071],prg0[1069],prg0[1067],prg0[1065],prg0[1063],prg0[1061],prg0[1059],prg0[1057],
                prg0[1070],prg0[1068],prg0[1066],prg0[1064],prg0[1062],prg0[1060],prg0[1058],prg0[1056],
                prg0[1055],prg0[1053],prg0[1051],prg0[1049],prg0[1047],prg0[1045],prg0[1043],prg0[1041],
                prg0[1054],prg0[1052],prg0[1050],prg0[1048],prg0[1046],prg0[1044],prg0[1042],prg0[1040],
                prg0[1039],prg0[1037],prg0[1035],prg0[1033],prg0[1031],prg0[1029],prg0[1027],prg0[1025],
                prg0[1038],prg0[1036],prg0[1034],prg0[1032],prg0[1030],prg0[1028],prg0[1026],prg0[1024]}),
       .INIT_3({prg0[1023],prg0[1021],prg0[1019],prg0[1017],prg0[1015],prg0[1013],prg0[1011],prg0[1009],
                prg0[1022],prg0[1020],prg0[1018],prg0[1016],prg0[1014],prg0[1012],prg0[1010],prg0[1008],
                prg0[1007],prg0[1005],prg0[1003],prg0[1001],prg0[ 999],prg0[ 997],prg0[ 995],prg0[ 993],
                prg0[1006],prg0[1004],prg0[1002],prg0[1000],prg0[ 998],prg0[ 996],prg0[ 994],prg0[ 992],
                prg0[ 991],prg0[ 989],prg0[ 987],prg0[ 985],prg0[ 983],prg0[ 981],prg0[ 979],prg0[ 977],
                prg0[ 990],prg0[ 988],prg0[ 986],prg0[ 984],prg0[ 982],prg0[ 980],prg0[ 978],prg0[ 976],
                prg0[ 975],prg0[ 973],prg0[ 971],prg0[ 969],prg0[ 967],prg0[ 965],prg0[ 963],prg0[ 961],
                prg0[ 974],prg0[ 972],prg0[ 970],prg0[ 968],prg0[ 966],prg0[ 964],prg0[ 962],prg0[ 960],
                prg0[ 959],prg0[ 957],prg0[ 955],prg0[ 953],prg0[ 951],prg0[ 949],prg0[ 947],prg0[ 945],
                prg0[ 958],prg0[ 956],prg0[ 954],prg0[ 952],prg0[ 950],prg0[ 948],prg0[ 946],prg0[ 944],
                prg0[ 943],prg0[ 941],prg0[ 939],prg0[ 937],prg0[ 935],prg0[ 933],prg0[ 931],prg0[ 929],
                prg0[ 942],prg0[ 940],prg0[ 938],prg0[ 936],prg0[ 934],prg0[ 932],prg0[ 930],prg0[ 928],
                prg0[ 927],prg0[ 925],prg0[ 923],prg0[ 921],prg0[ 919],prg0[ 917],prg0[ 915],prg0[ 913],
                prg0[ 926],prg0[ 924],prg0[ 922],prg0[ 920],prg0[ 918],prg0[ 916],prg0[ 914],prg0[ 912],
                prg0[ 911],prg0[ 909],prg0[ 907],prg0[ 905],prg0[ 903],prg0[ 901],prg0[ 899],prg0[ 897],
                prg0[ 910],prg0[ 908],prg0[ 906],prg0[ 904],prg0[ 902],prg0[ 900],prg0[ 898],prg0[ 896],
                prg0[ 895],prg0[ 893],prg0[ 891],prg0[ 889],prg0[ 887],prg0[ 885],prg0[ 883],prg0[ 881],
                prg0[ 894],prg0[ 892],prg0[ 890],prg0[ 888],prg0[ 886],prg0[ 884],prg0[ 882],prg0[ 880],
                prg0[ 879],prg0[ 877],prg0[ 875],prg0[ 873],prg0[ 871],prg0[ 869],prg0[ 867],prg0[ 865],
                prg0[ 878],prg0[ 876],prg0[ 874],prg0[ 872],prg0[ 870],prg0[ 868],prg0[ 866],prg0[ 864],
                prg0[ 863],prg0[ 861],prg0[ 859],prg0[ 857],prg0[ 855],prg0[ 853],prg0[ 851],prg0[ 849],
                prg0[ 862],prg0[ 860],prg0[ 858],prg0[ 856],prg0[ 854],prg0[ 852],prg0[ 850],prg0[ 848],
                prg0[ 847],prg0[ 845],prg0[ 843],prg0[ 841],prg0[ 839],prg0[ 837],prg0[ 835],prg0[ 833],
                prg0[ 846],prg0[ 844],prg0[ 842],prg0[ 840],prg0[ 838],prg0[ 836],prg0[ 834],prg0[ 832],
                prg0[ 831],prg0[ 829],prg0[ 827],prg0[ 825],prg0[ 823],prg0[ 821],prg0[ 819],prg0[ 817],
                prg0[ 830],prg0[ 828],prg0[ 826],prg0[ 824],prg0[ 822],prg0[ 820],prg0[ 818],prg0[ 816],
                prg0[ 815],prg0[ 813],prg0[ 811],prg0[ 809],prg0[ 807],prg0[ 805],prg0[ 803],prg0[ 801],
                prg0[ 814],prg0[ 812],prg0[ 810],prg0[ 808],prg0[ 806],prg0[ 804],prg0[ 802],prg0[ 800],
                prg0[ 799],prg0[ 797],prg0[ 795],prg0[ 793],prg0[ 791],prg0[ 789],prg0[ 787],prg0[ 785],
                prg0[ 798],prg0[ 796],prg0[ 794],prg0[ 792],prg0[ 790],prg0[ 788],prg0[ 786],prg0[ 784],
                prg0[ 783],prg0[ 781],prg0[ 779],prg0[ 777],prg0[ 775],prg0[ 773],prg0[ 771],prg0[ 769],
                prg0[ 782],prg0[ 780],prg0[ 778],prg0[ 776],prg0[ 774],prg0[ 772],prg0[ 770],prg0[ 768]}),
       .INIT_2({prg0[ 767],prg0[ 765],prg0[ 763],prg0[ 761],prg0[ 759],prg0[ 757],prg0[ 755],prg0[ 753],
                prg0[ 766],prg0[ 764],prg0[ 762],prg0[ 760],prg0[ 758],prg0[ 756],prg0[ 754],prg0[ 752],
                prg0[ 751],prg0[ 749],prg0[ 747],prg0[ 745],prg0[ 743],prg0[ 741],prg0[ 739],prg0[ 737],
                prg0[ 750],prg0[ 748],prg0[ 746],prg0[ 744],prg0[ 742],prg0[ 740],prg0[ 738],prg0[ 736],
                prg0[ 735],prg0[ 733],prg0[ 731],prg0[ 729],prg0[ 727],prg0[ 725],prg0[ 723],prg0[ 721],
                prg0[ 734],prg0[ 732],prg0[ 730],prg0[ 728],prg0[ 726],prg0[ 724],prg0[ 722],prg0[ 720],
                prg0[ 719],prg0[ 717],prg0[ 715],prg0[ 713],prg0[ 711],prg0[ 709],prg0[ 707],prg0[ 705],
                prg0[ 718],prg0[ 716],prg0[ 714],prg0[ 712],prg0[ 710],prg0[ 708],prg0[ 706],prg0[ 704],
                prg0[ 703],prg0[ 701],prg0[ 699],prg0[ 697],prg0[ 695],prg0[ 693],prg0[ 691],prg0[ 689],
                prg0[ 702],prg0[ 700],prg0[ 698],prg0[ 696],prg0[ 694],prg0[ 692],prg0[ 690],prg0[ 688],
                prg0[ 687],prg0[ 685],prg0[ 683],prg0[ 681],prg0[ 679],prg0[ 677],prg0[ 675],prg0[ 673],
                prg0[ 686],prg0[ 684],prg0[ 682],prg0[ 680],prg0[ 678],prg0[ 676],prg0[ 674],prg0[ 672],
                prg0[ 671],prg0[ 669],prg0[ 667],prg0[ 665],prg0[ 663],prg0[ 661],prg0[ 659],prg0[ 657],
                prg0[ 670],prg0[ 668],prg0[ 666],prg0[ 664],prg0[ 662],prg0[ 660],prg0[ 658],prg0[ 656],
                prg0[ 655],prg0[ 653],prg0[ 651],prg0[ 649],prg0[ 647],prg0[ 645],prg0[ 643],prg0[ 641],
                prg0[ 654],prg0[ 652],prg0[ 650],prg0[ 648],prg0[ 646],prg0[ 644],prg0[ 642],prg0[ 640],
                prg0[ 639],prg0[ 637],prg0[ 635],prg0[ 633],prg0[ 631],prg0[ 629],prg0[ 627],prg0[ 625],
                prg0[ 638],prg0[ 636],prg0[ 634],prg0[ 632],prg0[ 630],prg0[ 628],prg0[ 626],prg0[ 624],
                prg0[ 623],prg0[ 621],prg0[ 619],prg0[ 617],prg0[ 615],prg0[ 613],prg0[ 611],prg0[ 609],
                prg0[ 622],prg0[ 620],prg0[ 618],prg0[ 616],prg0[ 614],prg0[ 612],prg0[ 610],prg0[ 608],
                prg0[ 607],prg0[ 605],prg0[ 603],prg0[ 601],prg0[ 599],prg0[ 597],prg0[ 595],prg0[ 593],
                prg0[ 606],prg0[ 604],prg0[ 602],prg0[ 600],prg0[ 598],prg0[ 596],prg0[ 594],prg0[ 592],
                prg0[ 591],prg0[ 589],prg0[ 587],prg0[ 585],prg0[ 583],prg0[ 581],prg0[ 579],prg0[ 577],
                prg0[ 590],prg0[ 588],prg0[ 586],prg0[ 584],prg0[ 582],prg0[ 580],prg0[ 578],prg0[ 576],
                prg0[ 575],prg0[ 573],prg0[ 571],prg0[ 569],prg0[ 567],prg0[ 565],prg0[ 563],prg0[ 561],
                prg0[ 574],prg0[ 572],prg0[ 570],prg0[ 568],prg0[ 566],prg0[ 564],prg0[ 562],prg0[ 560],
                prg0[ 559],prg0[ 557],prg0[ 555],prg0[ 553],prg0[ 551],prg0[ 549],prg0[ 547],prg0[ 545],
                prg0[ 558],prg0[ 556],prg0[ 554],prg0[ 552],prg0[ 550],prg0[ 548],prg0[ 546],prg0[ 544],
                prg0[ 543],prg0[ 541],prg0[ 539],prg0[ 537],prg0[ 535],prg0[ 533],prg0[ 531],prg0[ 529],
                prg0[ 542],prg0[ 540],prg0[ 538],prg0[ 536],prg0[ 534],prg0[ 532],prg0[ 530],prg0[ 528],
                prg0[ 527],prg0[ 525],prg0[ 523],prg0[ 521],prg0[ 519],prg0[ 517],prg0[ 515],prg0[ 513],
                prg0[ 526],prg0[ 524],prg0[ 522],prg0[ 520],prg0[ 518],prg0[ 516],prg0[ 514],prg0[ 512]}),
       .INIT_1({prg0[ 511],prg0[ 509],prg0[ 507],prg0[ 505],prg0[ 503],prg0[ 501],prg0[ 499],prg0[ 497],
                prg0[ 510],prg0[ 508],prg0[ 506],prg0[ 504],prg0[ 502],prg0[ 500],prg0[ 498],prg0[ 496],
                prg0[ 495],prg0[ 493],prg0[ 491],prg0[ 489],prg0[ 487],prg0[ 485],prg0[ 483],prg0[ 481],
                prg0[ 494],prg0[ 492],prg0[ 490],prg0[ 488],prg0[ 486],prg0[ 484],prg0[ 482],prg0[ 480],
                prg0[ 479],prg0[ 477],prg0[ 475],prg0[ 473],prg0[ 471],prg0[ 469],prg0[ 467],prg0[ 465],
                prg0[ 478],prg0[ 476],prg0[ 474],prg0[ 472],prg0[ 470],prg0[ 468],prg0[ 466],prg0[ 464],
                prg0[ 463],prg0[ 461],prg0[ 459],prg0[ 457],prg0[ 455],prg0[ 453],prg0[ 451],prg0[ 449],
                prg0[ 462],prg0[ 460],prg0[ 458],prg0[ 456],prg0[ 454],prg0[ 452],prg0[ 450],prg0[ 448],
                prg0[ 447],prg0[ 445],prg0[ 443],prg0[ 441],prg0[ 439],prg0[ 437],prg0[ 435],prg0[ 433],
                prg0[ 446],prg0[ 444],prg0[ 442],prg0[ 440],prg0[ 438],prg0[ 436],prg0[ 434],prg0[ 432],
                prg0[ 431],prg0[ 429],prg0[ 427],prg0[ 425],prg0[ 423],prg0[ 421],prg0[ 419],prg0[ 417],
                prg0[ 430],prg0[ 428],prg0[ 426],prg0[ 424],prg0[ 422],prg0[ 420],prg0[ 418],prg0[ 416],
                prg0[ 415],prg0[ 413],prg0[ 411],prg0[ 409],prg0[ 407],prg0[ 405],prg0[ 403],prg0[ 401],
                prg0[ 414],prg0[ 412],prg0[ 410],prg0[ 408],prg0[ 406],prg0[ 404],prg0[ 402],prg0[ 400],
                prg0[ 399],prg0[ 397],prg0[ 395],prg0[ 393],prg0[ 391],prg0[ 389],prg0[ 387],prg0[ 385],
                prg0[ 398],prg0[ 396],prg0[ 394],prg0[ 392],prg0[ 390],prg0[ 388],prg0[ 386],prg0[ 384],
                prg0[ 383],prg0[ 381],prg0[ 379],prg0[ 377],prg0[ 375],prg0[ 373],prg0[ 371],prg0[ 369],
                prg0[ 382],prg0[ 380],prg0[ 378],prg0[ 376],prg0[ 374],prg0[ 372],prg0[ 370],prg0[ 368],
                prg0[ 367],prg0[ 365],prg0[ 363],prg0[ 361],prg0[ 359],prg0[ 357],prg0[ 355],prg0[ 353],
                prg0[ 366],prg0[ 364],prg0[ 362],prg0[ 360],prg0[ 358],prg0[ 356],prg0[ 354],prg0[ 352],
                prg0[ 351],prg0[ 349],prg0[ 347],prg0[ 345],prg0[ 343],prg0[ 341],prg0[ 339],prg0[ 337],
                prg0[ 350],prg0[ 348],prg0[ 346],prg0[ 344],prg0[ 342],prg0[ 340],prg0[ 338],prg0[ 336],
                prg0[ 335],prg0[ 333],prg0[ 331],prg0[ 329],prg0[ 327],prg0[ 325],prg0[ 323],prg0[ 321],
                prg0[ 334],prg0[ 332],prg0[ 330],prg0[ 328],prg0[ 326],prg0[ 324],prg0[ 322],prg0[ 320],
                prg0[ 319],prg0[ 317],prg0[ 315],prg0[ 313],prg0[ 311],prg0[ 309],prg0[ 307],prg0[ 305],
                prg0[ 318],prg0[ 316],prg0[ 314],prg0[ 312],prg0[ 310],prg0[ 308],prg0[ 306],prg0[ 304],
                prg0[ 303],prg0[ 301],prg0[ 299],prg0[ 297],prg0[ 295],prg0[ 293],prg0[ 291],prg0[ 289],
                prg0[ 302],prg0[ 300],prg0[ 298],prg0[ 296],prg0[ 294],prg0[ 292],prg0[ 290],prg0[ 288],
                prg0[ 287],prg0[ 285],prg0[ 283],prg0[ 281],prg0[ 279],prg0[ 277],prg0[ 275],prg0[ 273],
                prg0[ 286],prg0[ 284],prg0[ 282],prg0[ 280],prg0[ 278],prg0[ 276],prg0[ 274],prg0[ 272],
                prg0[ 271],prg0[ 269],prg0[ 267],prg0[ 265],prg0[ 263],prg0[ 261],prg0[ 259],prg0[ 257],
                prg0[ 270],prg0[ 268],prg0[ 266],prg0[ 264],prg0[ 262],prg0[ 260],prg0[ 258],prg0[ 256]}),
       .INIT_0({prg0[ 255],prg0[ 253],prg0[ 251],prg0[ 249],prg0[ 247],prg0[ 245],prg0[ 243],prg0[ 241],
                prg0[ 254],prg0[ 252],prg0[ 250],prg0[ 248],prg0[ 246],prg0[ 244],prg0[ 242],prg0[ 240],
                prg0[ 239],prg0[ 237],prg0[ 235],prg0[ 233],prg0[ 231],prg0[ 229],prg0[ 227],prg0[ 225],
                prg0[ 238],prg0[ 236],prg0[ 234],prg0[ 232],prg0[ 230],prg0[ 228],prg0[ 226],prg0[ 224],
                prg0[ 223],prg0[ 221],prg0[ 219],prg0[ 217],prg0[ 215],prg0[ 213],prg0[ 211],prg0[ 209],
                prg0[ 222],prg0[ 220],prg0[ 218],prg0[ 216],prg0[ 214],prg0[ 212],prg0[ 210],prg0[ 208],
                prg0[ 207],prg0[ 205],prg0[ 203],prg0[ 201],prg0[ 199],prg0[ 197],prg0[ 195],prg0[ 193],
                prg0[ 206],prg0[ 204],prg0[ 202],prg0[ 200],prg0[ 198],prg0[ 196],prg0[ 194],prg0[ 192],
                prg0[ 191],prg0[ 189],prg0[ 187],prg0[ 185],prg0[ 183],prg0[ 181],prg0[ 179],prg0[ 177],
                prg0[ 190],prg0[ 188],prg0[ 186],prg0[ 184],prg0[ 182],prg0[ 180],prg0[ 178],prg0[ 176],
                prg0[ 175],prg0[ 173],prg0[ 171],prg0[ 169],prg0[ 167],prg0[ 165],prg0[ 163],prg0[ 161],
                prg0[ 174],prg0[ 172],prg0[ 170],prg0[ 168],prg0[ 166],prg0[ 164],prg0[ 162],prg0[ 160],
                prg0[ 159],prg0[ 157],prg0[ 155],prg0[ 153],prg0[ 151],prg0[ 149],prg0[ 147],prg0[ 145],
                prg0[ 158],prg0[ 156],prg0[ 154],prg0[ 152],prg0[ 150],prg0[ 148],prg0[ 146],prg0[ 144],
                prg0[ 143],prg0[ 141],prg0[ 139],prg0[ 137],prg0[ 135],prg0[ 133],prg0[ 131],prg0[ 129],
                prg0[ 142],prg0[ 140],prg0[ 138],prg0[ 136],prg0[ 134],prg0[ 132],prg0[ 130],prg0[ 128],
                prg0[ 127],prg0[ 125],prg0[ 123],prg0[ 121],prg0[ 119],prg0[ 117],prg0[ 115],prg0[ 113],
                prg0[ 126],prg0[ 124],prg0[ 122],prg0[ 120],prg0[ 118],prg0[ 116],prg0[ 114],prg0[ 112],
                prg0[ 111],prg0[ 109],prg0[ 107],prg0[ 105],prg0[ 103],prg0[ 101],prg0[  99],prg0[  97],
                prg0[ 110],prg0[ 108],prg0[ 106],prg0[ 104],prg0[ 102],prg0[ 100],prg0[  98],prg0[  96],
                prg0[  95],prg0[  93],prg0[  91],prg0[  89],prg0[  87],prg0[  85],prg0[  83],prg0[  81],
                prg0[  94],prg0[  92],prg0[  90],prg0[  88],prg0[  86],prg0[  84],prg0[  82],prg0[  80],
                prg0[  79],prg0[  77],prg0[  75],prg0[  73],prg0[  71],prg0[  69],prg0[  67],prg0[  65],
                prg0[  78],prg0[  76],prg0[  74],prg0[  72],prg0[  70],prg0[  68],prg0[  66],prg0[  64],
                prg0[  63],prg0[  61],prg0[  59],prg0[  57],prg0[  55],prg0[  53],prg0[  51],prg0[  49],
                prg0[  62],prg0[  60],prg0[  58],prg0[  56],prg0[  54],prg0[  52],prg0[  50],prg0[  48],
                prg0[  47],prg0[  45],prg0[  43],prg0[  41],prg0[  39],prg0[  37],prg0[  35],prg0[  33],
                prg0[  46],prg0[  44],prg0[  42],prg0[  40],prg0[  38],prg0[  36],prg0[  34],prg0[  32],
                prg0[  31],prg0[  29],prg0[  27],prg0[  25],prg0[  23],prg0[  21],prg0[  19],prg0[  17],
                prg0[  30],prg0[  28],prg0[  26],prg0[  24],prg0[  22],prg0[  20],prg0[  18],prg0[  16],
                prg0[  15],prg0[  13],prg0[  11],prg0[   9],prg0[   7],prg0[   5],prg0[   3],prg0[   1],
                prg0[  14],prg0[  12],prg0[  10],prg0[   8],prg0[   6],prg0[   4],prg0[   2],prg0[   0]}),
       .READ_MODE(3),
       .WRITE_MODE(3))
   mem
     (// Outputs
      .RDATA  ( {dum14[13:10],
                 DAT_O[1],dum14[9:3],
                 DAT_O[0],dum14[2:0]}         ),
      // Input
      .MASK   ( 16'h0                         ),
      .WDATA  ( {4'h0,                       
                 B[1],7'h0,
                 B[0],3'b0}       ),                       
      .WADDR  ( {Wai[2:0],Wai[10:3]}          ), // Note mangling
      .RADDR  ( {Rai[2:0],Rai[10:3]}          ), // Note mangling
      .RE     ( 1'b1                          ),
      .WE     ( we                            ), 
      .WCLK   ( clk                           ),
      .RCLK   ( clk                           ),
      .RCLKE  ( 1'b1                          ),
      .WCLKE  ( 1'b1                          ) 
      /*AUTOINST*/);
   
endmodule
