/* -----------------------------------------------------------------------------
 * Part of midgetv
 * 2019. Copyright B. Nossum.
 * For licence, see LICENCE
 * -----------------------------------------------------------------------------
 * EBR program memory is split into 8-bit wide memory specified here.
 */
module m_ebr_w8
  # ( parameter EBRADRWIDTH = 9,
      parameter [4095:0] prg0 = 4096'h0,
      parameter [4095:0] prg1 = 4096'h0,
      parameter [4095:0] prg2 = 4096'h0,
      parameter [4095:0] prg3 = 4096'h0
      )
   (
    input [7:0]             B, //     Output from ALU
    input [EBRADRWIDTH-1:0] Rai, //   Read address
    input [EBRADRWIDTH-1:0] Wai, //   Write address
    input                   clk, //   System clock
    input                   bmask, // Byte mask for write, active LUW
    input                   iwe, //   Write enable
    output [7:0]            DAT_O //  Registered output
    );
   wire                     we = ~bmask & iwe;
   
   localparam NrRamsHere = (1<<(EBRADRWIDTH-9));

   generate

      if ( NrRamsHere == 1 ) begin
         /* verilator lint_off UNUSED */
         wire [7:0] dum8;
         /* verilator lint_on UNUSED */

         SB_RAM40_4K 
           #(
             .INIT_F({prg0[4095],prg0[4087],prg0[4094],prg0[4086],prg0[4093],prg0[4085],prg0[4092],prg0[4084],
                      prg0[4091],prg0[4083],prg0[4090],prg0[4082],prg0[4089],prg0[4081],prg0[4088],prg0[4080],
                      prg0[4079],prg0[4071],prg0[4078],prg0[4070],prg0[4077],prg0[4069],prg0[4076],prg0[4068],
                      prg0[4075],prg0[4067],prg0[4074],prg0[4066],prg0[4073],prg0[4065],prg0[4072],prg0[4064],
                      prg0[4063],prg0[4055],prg0[4062],prg0[4054],prg0[4061],prg0[4053],prg0[4060],prg0[4052],
                      prg0[4059],prg0[4051],prg0[4058],prg0[4050],prg0[4057],prg0[4049],prg0[4056],prg0[4048],
                      prg0[4047],prg0[4039],prg0[4046],prg0[4038],prg0[4045],prg0[4037],prg0[4044],prg0[4036],
                      prg0[4043],prg0[4035],prg0[4042],prg0[4034],prg0[4041],prg0[4033],prg0[4040],prg0[4032],
                      prg0[4031],prg0[4023],prg0[4030],prg0[4022],prg0[4029],prg0[4021],prg0[4028],prg0[4020],
                      prg0[4027],prg0[4019],prg0[4026],prg0[4018],prg0[4025],prg0[4017],prg0[4024],prg0[4016],
                      prg0[4015],prg0[4007],prg0[4014],prg0[4006],prg0[4013],prg0[4005],prg0[4012],prg0[4004],
                      prg0[4011],prg0[4003],prg0[4010],prg0[4002],prg0[4009],prg0[4001],prg0[4008],prg0[4000],
                      prg0[3999],prg0[3991],prg0[3998],prg0[3990],prg0[3997],prg0[3989],prg0[3996],prg0[3988],
                      prg0[3995],prg0[3987],prg0[3994],prg0[3986],prg0[3993],prg0[3985],prg0[3992],prg0[3984],
                      prg0[3983],prg0[3975],prg0[3982],prg0[3974],prg0[3981],prg0[3973],prg0[3980],prg0[3972],
                      prg0[3979],prg0[3971],prg0[3978],prg0[3970],prg0[3977],prg0[3969],prg0[3976],prg0[3968],
                      prg0[3967],prg0[3959],prg0[3966],prg0[3958],prg0[3965],prg0[3957],prg0[3964],prg0[3956],
                      prg0[3963],prg0[3955],prg0[3962],prg0[3954],prg0[3961],prg0[3953],prg0[3960],prg0[3952],
                      prg0[3951],prg0[3943],prg0[3950],prg0[3942],prg0[3949],prg0[3941],prg0[3948],prg0[3940],
                      prg0[3947],prg0[3939],prg0[3946],prg0[3938],prg0[3945],prg0[3937],prg0[3944],prg0[3936],
                      prg0[3935],prg0[3927],prg0[3934],prg0[3926],prg0[3933],prg0[3925],prg0[3932],prg0[3924],
                      prg0[3931],prg0[3923],prg0[3930],prg0[3922],prg0[3929],prg0[3921],prg0[3928],prg0[3920],
                      prg0[3919],prg0[3911],prg0[3918],prg0[3910],prg0[3917],prg0[3909],prg0[3916],prg0[3908],
                      prg0[3915],prg0[3907],prg0[3914],prg0[3906],prg0[3913],prg0[3905],prg0[3912],prg0[3904],
                      prg0[3903],prg0[3895],prg0[3902],prg0[3894],prg0[3901],prg0[3893],prg0[3900],prg0[3892],
                      prg0[3899],prg0[3891],prg0[3898],prg0[3890],prg0[3897],prg0[3889],prg0[3896],prg0[3888],
                      prg0[3887],prg0[3879],prg0[3886],prg0[3878],prg0[3885],prg0[3877],prg0[3884],prg0[3876],
                      prg0[3883],prg0[3875],prg0[3882],prg0[3874],prg0[3881],prg0[3873],prg0[3880],prg0[3872],
                      prg0[3871],prg0[3863],prg0[3870],prg0[3862],prg0[3869],prg0[3861],prg0[3868],prg0[3860],
                      prg0[3867],prg0[3859],prg0[3866],prg0[3858],prg0[3865],prg0[3857],prg0[3864],prg0[3856],
                      prg0[3855],prg0[3847],prg0[3854],prg0[3846],prg0[3853],prg0[3845],prg0[3852],prg0[3844],
                      prg0[3851],prg0[3843],prg0[3850],prg0[3842],prg0[3849],prg0[3841],prg0[3848],prg0[3840]}),
             .INIT_E({prg0[3839],prg0[3831],prg0[3838],prg0[3830],prg0[3837],prg0[3829],prg0[3836],prg0[3828],
                      prg0[3835],prg0[3827],prg0[3834],prg0[3826],prg0[3833],prg0[3825],prg0[3832],prg0[3824],
                      prg0[3823],prg0[3815],prg0[3822],prg0[3814],prg0[3821],prg0[3813],prg0[3820],prg0[3812],
                      prg0[3819],prg0[3811],prg0[3818],prg0[3810],prg0[3817],prg0[3809],prg0[3816],prg0[3808],
                      prg0[3807],prg0[3799],prg0[3806],prg0[3798],prg0[3805],prg0[3797],prg0[3804],prg0[3796],
                      prg0[3803],prg0[3795],prg0[3802],prg0[3794],prg0[3801],prg0[3793],prg0[3800],prg0[3792],
                      prg0[3791],prg0[3783],prg0[3790],prg0[3782],prg0[3789],prg0[3781],prg0[3788],prg0[3780],
                      prg0[3787],prg0[3779],prg0[3786],prg0[3778],prg0[3785],prg0[3777],prg0[3784],prg0[3776],
                      prg0[3775],prg0[3767],prg0[3774],prg0[3766],prg0[3773],prg0[3765],prg0[3772],prg0[3764],
                      prg0[3771],prg0[3763],prg0[3770],prg0[3762],prg0[3769],prg0[3761],prg0[3768],prg0[3760],
                      prg0[3759],prg0[3751],prg0[3758],prg0[3750],prg0[3757],prg0[3749],prg0[3756],prg0[3748],
                      prg0[3755],prg0[3747],prg0[3754],prg0[3746],prg0[3753],prg0[3745],prg0[3752],prg0[3744],
                      prg0[3743],prg0[3735],prg0[3742],prg0[3734],prg0[3741],prg0[3733],prg0[3740],prg0[3732],
                      prg0[3739],prg0[3731],prg0[3738],prg0[3730],prg0[3737],prg0[3729],prg0[3736],prg0[3728],
                      prg0[3727],prg0[3719],prg0[3726],prg0[3718],prg0[3725],prg0[3717],prg0[3724],prg0[3716],
                      prg0[3723],prg0[3715],prg0[3722],prg0[3714],prg0[3721],prg0[3713],prg0[3720],prg0[3712],
                      prg0[3711],prg0[3703],prg0[3710],prg0[3702],prg0[3709],prg0[3701],prg0[3708],prg0[3700],
                      prg0[3707],prg0[3699],prg0[3706],prg0[3698],prg0[3705],prg0[3697],prg0[3704],prg0[3696],
                      prg0[3695],prg0[3687],prg0[3694],prg0[3686],prg0[3693],prg0[3685],prg0[3692],prg0[3684],
                      prg0[3691],prg0[3683],prg0[3690],prg0[3682],prg0[3689],prg0[3681],prg0[3688],prg0[3680],
                      prg0[3679],prg0[3671],prg0[3678],prg0[3670],prg0[3677],prg0[3669],prg0[3676],prg0[3668],
                      prg0[3675],prg0[3667],prg0[3674],prg0[3666],prg0[3673],prg0[3665],prg0[3672],prg0[3664],
                      prg0[3663],prg0[3655],prg0[3662],prg0[3654],prg0[3661],prg0[3653],prg0[3660],prg0[3652],
                      prg0[3659],prg0[3651],prg0[3658],prg0[3650],prg0[3657],prg0[3649],prg0[3656],prg0[3648],
                      prg0[3647],prg0[3639],prg0[3646],prg0[3638],prg0[3645],prg0[3637],prg0[3644],prg0[3636],
                      prg0[3643],prg0[3635],prg0[3642],prg0[3634],prg0[3641],prg0[3633],prg0[3640],prg0[3632],
                      prg0[3631],prg0[3623],prg0[3630],prg0[3622],prg0[3629],prg0[3621],prg0[3628],prg0[3620],
                      prg0[3627],prg0[3619],prg0[3626],prg0[3618],prg0[3625],prg0[3617],prg0[3624],prg0[3616],
                      prg0[3615],prg0[3607],prg0[3614],prg0[3606],prg0[3613],prg0[3605],prg0[3612],prg0[3604],
                      prg0[3611],prg0[3603],prg0[3610],prg0[3602],prg0[3609],prg0[3601],prg0[3608],prg0[3600],
                      prg0[3599],prg0[3591],prg0[3598],prg0[3590],prg0[3597],prg0[3589],prg0[3596],prg0[3588],
                      prg0[3595],prg0[3587],prg0[3594],prg0[3586],prg0[3593],prg0[3585],prg0[3592],prg0[3584]}),
             .INIT_D({prg0[3583],prg0[3575],prg0[3582],prg0[3574],prg0[3581],prg0[3573],prg0[3580],prg0[3572],
                      prg0[3579],prg0[3571],prg0[3578],prg0[3570],prg0[3577],prg0[3569],prg0[3576],prg0[3568],
                      prg0[3567],prg0[3559],prg0[3566],prg0[3558],prg0[3565],prg0[3557],prg0[3564],prg0[3556],
                      prg0[3563],prg0[3555],prg0[3562],prg0[3554],prg0[3561],prg0[3553],prg0[3560],prg0[3552],
                      prg0[3551],prg0[3543],prg0[3550],prg0[3542],prg0[3549],prg0[3541],prg0[3548],prg0[3540],
                      prg0[3547],prg0[3539],prg0[3546],prg0[3538],prg0[3545],prg0[3537],prg0[3544],prg0[3536],
                      prg0[3535],prg0[3527],prg0[3534],prg0[3526],prg0[3533],prg0[3525],prg0[3532],prg0[3524],
                      prg0[3531],prg0[3523],prg0[3530],prg0[3522],prg0[3529],prg0[3521],prg0[3528],prg0[3520],
                      prg0[3519],prg0[3511],prg0[3518],prg0[3510],prg0[3517],prg0[3509],prg0[3516],prg0[3508],
                      prg0[3515],prg0[3507],prg0[3514],prg0[3506],prg0[3513],prg0[3505],prg0[3512],prg0[3504],
                      prg0[3503],prg0[3495],prg0[3502],prg0[3494],prg0[3501],prg0[3493],prg0[3500],prg0[3492],
                      prg0[3499],prg0[3491],prg0[3498],prg0[3490],prg0[3497],prg0[3489],prg0[3496],prg0[3488],
                      prg0[3487],prg0[3479],prg0[3486],prg0[3478],prg0[3485],prg0[3477],prg0[3484],prg0[3476],
                      prg0[3483],prg0[3475],prg0[3482],prg0[3474],prg0[3481],prg0[3473],prg0[3480],prg0[3472],
                      prg0[3471],prg0[3463],prg0[3470],prg0[3462],prg0[3469],prg0[3461],prg0[3468],prg0[3460],
                      prg0[3467],prg0[3459],prg0[3466],prg0[3458],prg0[3465],prg0[3457],prg0[3464],prg0[3456],
                      prg0[3455],prg0[3447],prg0[3454],prg0[3446],prg0[3453],prg0[3445],prg0[3452],prg0[3444],
                      prg0[3451],prg0[3443],prg0[3450],prg0[3442],prg0[3449],prg0[3441],prg0[3448],prg0[3440],
                      prg0[3439],prg0[3431],prg0[3438],prg0[3430],prg0[3437],prg0[3429],prg0[3436],prg0[3428],
                      prg0[3435],prg0[3427],prg0[3434],prg0[3426],prg0[3433],prg0[3425],prg0[3432],prg0[3424],
                      prg0[3423],prg0[3415],prg0[3422],prg0[3414],prg0[3421],prg0[3413],prg0[3420],prg0[3412],
                      prg0[3419],prg0[3411],prg0[3418],prg0[3410],prg0[3417],prg0[3409],prg0[3416],prg0[3408],
                      prg0[3407],prg0[3399],prg0[3406],prg0[3398],prg0[3405],prg0[3397],prg0[3404],prg0[3396],
                      prg0[3403],prg0[3395],prg0[3402],prg0[3394],prg0[3401],prg0[3393],prg0[3400],prg0[3392],
                      prg0[3391],prg0[3383],prg0[3390],prg0[3382],prg0[3389],prg0[3381],prg0[3388],prg0[3380],
                      prg0[3387],prg0[3379],prg0[3386],prg0[3378],prg0[3385],prg0[3377],prg0[3384],prg0[3376],
                      prg0[3375],prg0[3367],prg0[3374],prg0[3366],prg0[3373],prg0[3365],prg0[3372],prg0[3364],
                      prg0[3371],prg0[3363],prg0[3370],prg0[3362],prg0[3369],prg0[3361],prg0[3368],prg0[3360],
                      prg0[3359],prg0[3351],prg0[3358],prg0[3350],prg0[3357],prg0[3349],prg0[3356],prg0[3348],
                      prg0[3355],prg0[3347],prg0[3354],prg0[3346],prg0[3353],prg0[3345],prg0[3352],prg0[3344],
                      prg0[3343],prg0[3335],prg0[3342],prg0[3334],prg0[3341],prg0[3333],prg0[3340],prg0[3332],
                      prg0[3339],prg0[3331],prg0[3338],prg0[3330],prg0[3337],prg0[3329],prg0[3336],prg0[3328]}),
             .INIT_C({prg0[3327],prg0[3319],prg0[3326],prg0[3318],prg0[3325],prg0[3317],prg0[3324],prg0[3316],
                      prg0[3323],prg0[3315],prg0[3322],prg0[3314],prg0[3321],prg0[3313],prg0[3320],prg0[3312],
                      prg0[3311],prg0[3303],prg0[3310],prg0[3302],prg0[3309],prg0[3301],prg0[3308],prg0[3300],
                      prg0[3307],prg0[3299],prg0[3306],prg0[3298],prg0[3305],prg0[3297],prg0[3304],prg0[3296],
                      prg0[3295],prg0[3287],prg0[3294],prg0[3286],prg0[3293],prg0[3285],prg0[3292],prg0[3284],
                      prg0[3291],prg0[3283],prg0[3290],prg0[3282],prg0[3289],prg0[3281],prg0[3288],prg0[3280],
                      prg0[3279],prg0[3271],prg0[3278],prg0[3270],prg0[3277],prg0[3269],prg0[3276],prg0[3268],
                      prg0[3275],prg0[3267],prg0[3274],prg0[3266],prg0[3273],prg0[3265],prg0[3272],prg0[3264],
                      prg0[3263],prg0[3255],prg0[3262],prg0[3254],prg0[3261],prg0[3253],prg0[3260],prg0[3252],
                      prg0[3259],prg0[3251],prg0[3258],prg0[3250],prg0[3257],prg0[3249],prg0[3256],prg0[3248],
                      prg0[3247],prg0[3239],prg0[3246],prg0[3238],prg0[3245],prg0[3237],prg0[3244],prg0[3236],
                      prg0[3243],prg0[3235],prg0[3242],prg0[3234],prg0[3241],prg0[3233],prg0[3240],prg0[3232],
                      prg0[3231],prg0[3223],prg0[3230],prg0[3222],prg0[3229],prg0[3221],prg0[3228],prg0[3220],
                      prg0[3227],prg0[3219],prg0[3226],prg0[3218],prg0[3225],prg0[3217],prg0[3224],prg0[3216],
                      prg0[3215],prg0[3207],prg0[3214],prg0[3206],prg0[3213],prg0[3205],prg0[3212],prg0[3204],
                      prg0[3211],prg0[3203],prg0[3210],prg0[3202],prg0[3209],prg0[3201],prg0[3208],prg0[3200],
                      prg0[3199],prg0[3191],prg0[3198],prg0[3190],prg0[3197],prg0[3189],prg0[3196],prg0[3188],
                      prg0[3195],prg0[3187],prg0[3194],prg0[3186],prg0[3193],prg0[3185],prg0[3192],prg0[3184],
                      prg0[3183],prg0[3175],prg0[3182],prg0[3174],prg0[3181],prg0[3173],prg0[3180],prg0[3172],
                      prg0[3179],prg0[3171],prg0[3178],prg0[3170],prg0[3177],prg0[3169],prg0[3176],prg0[3168],
                      prg0[3167],prg0[3159],prg0[3166],prg0[3158],prg0[3165],prg0[3157],prg0[3164],prg0[3156],
                      prg0[3163],prg0[3155],prg0[3162],prg0[3154],prg0[3161],prg0[3153],prg0[3160],prg0[3152],
                      prg0[3151],prg0[3143],prg0[3150],prg0[3142],prg0[3149],prg0[3141],prg0[3148],prg0[3140],
                      prg0[3147],prg0[3139],prg0[3146],prg0[3138],prg0[3145],prg0[3137],prg0[3144],prg0[3136],
                      prg0[3135],prg0[3127],prg0[3134],prg0[3126],prg0[3133],prg0[3125],prg0[3132],prg0[3124],
                      prg0[3131],prg0[3123],prg0[3130],prg0[3122],prg0[3129],prg0[3121],prg0[3128],prg0[3120],
                      prg0[3119],prg0[3111],prg0[3118],prg0[3110],prg0[3117],prg0[3109],prg0[3116],prg0[3108],
                      prg0[3115],prg0[3107],prg0[3114],prg0[3106],prg0[3113],prg0[3105],prg0[3112],prg0[3104],
                      prg0[3103],prg0[3095],prg0[3102],prg0[3094],prg0[3101],prg0[3093],prg0[3100],prg0[3092],
                      prg0[3099],prg0[3091],prg0[3098],prg0[3090],prg0[3097],prg0[3089],prg0[3096],prg0[3088],
                      prg0[3087],prg0[3079],prg0[3086],prg0[3078],prg0[3085],prg0[3077],prg0[3084],prg0[3076],
                      prg0[3083],prg0[3075],prg0[3082],prg0[3074],prg0[3081],prg0[3073],prg0[3080],prg0[3072]}),
             .INIT_B({prg0[3071],prg0[3063],prg0[3070],prg0[3062],prg0[3069],prg0[3061],prg0[3068],prg0[3060],
                      prg0[3067],prg0[3059],prg0[3066],prg0[3058],prg0[3065],prg0[3057],prg0[3064],prg0[3056],
                      prg0[3055],prg0[3047],prg0[3054],prg0[3046],prg0[3053],prg0[3045],prg0[3052],prg0[3044],
                      prg0[3051],prg0[3043],prg0[3050],prg0[3042],prg0[3049],prg0[3041],prg0[3048],prg0[3040],
                      prg0[3039],prg0[3031],prg0[3038],prg0[3030],prg0[3037],prg0[3029],prg0[3036],prg0[3028],
                      prg0[3035],prg0[3027],prg0[3034],prg0[3026],prg0[3033],prg0[3025],prg0[3032],prg0[3024],
                      prg0[3023],prg0[3015],prg0[3022],prg0[3014],prg0[3021],prg0[3013],prg0[3020],prg0[3012],
                      prg0[3019],prg0[3011],prg0[3018],prg0[3010],prg0[3017],prg0[3009],prg0[3016],prg0[3008],
                      prg0[3007],prg0[2999],prg0[3006],prg0[2998],prg0[3005],prg0[2997],prg0[3004],prg0[2996],
                      prg0[3003],prg0[2995],prg0[3002],prg0[2994],prg0[3001],prg0[2993],prg0[3000],prg0[2992],
                      prg0[2991],prg0[2983],prg0[2990],prg0[2982],prg0[2989],prg0[2981],prg0[2988],prg0[2980],
                      prg0[2987],prg0[2979],prg0[2986],prg0[2978],prg0[2985],prg0[2977],prg0[2984],prg0[2976],
                      prg0[2975],prg0[2967],prg0[2974],prg0[2966],prg0[2973],prg0[2965],prg0[2972],prg0[2964],
                      prg0[2971],prg0[2963],prg0[2970],prg0[2962],prg0[2969],prg0[2961],prg0[2968],prg0[2960],
                      prg0[2959],prg0[2951],prg0[2958],prg0[2950],prg0[2957],prg0[2949],prg0[2956],prg0[2948],
                      prg0[2955],prg0[2947],prg0[2954],prg0[2946],prg0[2953],prg0[2945],prg0[2952],prg0[2944],
                      prg0[2943],prg0[2935],prg0[2942],prg0[2934],prg0[2941],prg0[2933],prg0[2940],prg0[2932],
                      prg0[2939],prg0[2931],prg0[2938],prg0[2930],prg0[2937],prg0[2929],prg0[2936],prg0[2928],
                      prg0[2927],prg0[2919],prg0[2926],prg0[2918],prg0[2925],prg0[2917],prg0[2924],prg0[2916],
                      prg0[2923],prg0[2915],prg0[2922],prg0[2914],prg0[2921],prg0[2913],prg0[2920],prg0[2912],
                      prg0[2911],prg0[2903],prg0[2910],prg0[2902],prg0[2909],prg0[2901],prg0[2908],prg0[2900],
                      prg0[2907],prg0[2899],prg0[2906],prg0[2898],prg0[2905],prg0[2897],prg0[2904],prg0[2896],
                      prg0[2895],prg0[2887],prg0[2894],prg0[2886],prg0[2893],prg0[2885],prg0[2892],prg0[2884],
                      prg0[2891],prg0[2883],prg0[2890],prg0[2882],prg0[2889],prg0[2881],prg0[2888],prg0[2880],
                      prg0[2879],prg0[2871],prg0[2878],prg0[2870],prg0[2877],prg0[2869],prg0[2876],prg0[2868],
                      prg0[2875],prg0[2867],prg0[2874],prg0[2866],prg0[2873],prg0[2865],prg0[2872],prg0[2864],
                      prg0[2863],prg0[2855],prg0[2862],prg0[2854],prg0[2861],prg0[2853],prg0[2860],prg0[2852],
                      prg0[2859],prg0[2851],prg0[2858],prg0[2850],prg0[2857],prg0[2849],prg0[2856],prg0[2848],
                      prg0[2847],prg0[2839],prg0[2846],prg0[2838],prg0[2845],prg0[2837],prg0[2844],prg0[2836],
                      prg0[2843],prg0[2835],prg0[2842],prg0[2834],prg0[2841],prg0[2833],prg0[2840],prg0[2832],
                      prg0[2831],prg0[2823],prg0[2830],prg0[2822],prg0[2829],prg0[2821],prg0[2828],prg0[2820],
                      prg0[2827],prg0[2819],prg0[2826],prg0[2818],prg0[2825],prg0[2817],prg0[2824],prg0[2816]}),
             .INIT_A({prg0[2815],prg0[2807],prg0[2814],prg0[2806],prg0[2813],prg0[2805],prg0[2812],prg0[2804],
                      prg0[2811],prg0[2803],prg0[2810],prg0[2802],prg0[2809],prg0[2801],prg0[2808],prg0[2800],
                      prg0[2799],prg0[2791],prg0[2798],prg0[2790],prg0[2797],prg0[2789],prg0[2796],prg0[2788],
                      prg0[2795],prg0[2787],prg0[2794],prg0[2786],prg0[2793],prg0[2785],prg0[2792],prg0[2784],
                      prg0[2783],prg0[2775],prg0[2782],prg0[2774],prg0[2781],prg0[2773],prg0[2780],prg0[2772],
                      prg0[2779],prg0[2771],prg0[2778],prg0[2770],prg0[2777],prg0[2769],prg0[2776],prg0[2768],
                      prg0[2767],prg0[2759],prg0[2766],prg0[2758],prg0[2765],prg0[2757],prg0[2764],prg0[2756],
                      prg0[2763],prg0[2755],prg0[2762],prg0[2754],prg0[2761],prg0[2753],prg0[2760],prg0[2752],
                      prg0[2751],prg0[2743],prg0[2750],prg0[2742],prg0[2749],prg0[2741],prg0[2748],prg0[2740],
                      prg0[2747],prg0[2739],prg0[2746],prg0[2738],prg0[2745],prg0[2737],prg0[2744],prg0[2736],
                      prg0[2735],prg0[2727],prg0[2734],prg0[2726],prg0[2733],prg0[2725],prg0[2732],prg0[2724],
                      prg0[2731],prg0[2723],prg0[2730],prg0[2722],prg0[2729],prg0[2721],prg0[2728],prg0[2720],
                      prg0[2719],prg0[2711],prg0[2718],prg0[2710],prg0[2717],prg0[2709],prg0[2716],prg0[2708],
                      prg0[2715],prg0[2707],prg0[2714],prg0[2706],prg0[2713],prg0[2705],prg0[2712],prg0[2704],
                      prg0[2703],prg0[2695],prg0[2702],prg0[2694],prg0[2701],prg0[2693],prg0[2700],prg0[2692],
                      prg0[2699],prg0[2691],prg0[2698],prg0[2690],prg0[2697],prg0[2689],prg0[2696],prg0[2688],
                      prg0[2687],prg0[2679],prg0[2686],prg0[2678],prg0[2685],prg0[2677],prg0[2684],prg0[2676],
                      prg0[2683],prg0[2675],prg0[2682],prg0[2674],prg0[2681],prg0[2673],prg0[2680],prg0[2672],
                      prg0[2671],prg0[2663],prg0[2670],prg0[2662],prg0[2669],prg0[2661],prg0[2668],prg0[2660],
                      prg0[2667],prg0[2659],prg0[2666],prg0[2658],prg0[2665],prg0[2657],prg0[2664],prg0[2656],
                      prg0[2655],prg0[2647],prg0[2654],prg0[2646],prg0[2653],prg0[2645],prg0[2652],prg0[2644],
                      prg0[2651],prg0[2643],prg0[2650],prg0[2642],prg0[2649],prg0[2641],prg0[2648],prg0[2640],
                      prg0[2639],prg0[2631],prg0[2638],prg0[2630],prg0[2637],prg0[2629],prg0[2636],prg0[2628],
                      prg0[2635],prg0[2627],prg0[2634],prg0[2626],prg0[2633],prg0[2625],prg0[2632],prg0[2624],
                      prg0[2623],prg0[2615],prg0[2622],prg0[2614],prg0[2621],prg0[2613],prg0[2620],prg0[2612],
                      prg0[2619],prg0[2611],prg0[2618],prg0[2610],prg0[2617],prg0[2609],prg0[2616],prg0[2608],
                      prg0[2607],prg0[2599],prg0[2606],prg0[2598],prg0[2605],prg0[2597],prg0[2604],prg0[2596],
                      prg0[2603],prg0[2595],prg0[2602],prg0[2594],prg0[2601],prg0[2593],prg0[2600],prg0[2592],
                      prg0[2591],prg0[2583],prg0[2590],prg0[2582],prg0[2589],prg0[2581],prg0[2588],prg0[2580],
                      prg0[2587],prg0[2579],prg0[2586],prg0[2578],prg0[2585],prg0[2577],prg0[2584],prg0[2576],
                      prg0[2575],prg0[2567],prg0[2574],prg0[2566],prg0[2573],prg0[2565],prg0[2572],prg0[2564],
                      prg0[2571],prg0[2563],prg0[2570],prg0[2562],prg0[2569],prg0[2561],prg0[2568],prg0[2560]}),
             .INIT_9({prg0[2559],prg0[2551],prg0[2558],prg0[2550],prg0[2557],prg0[2549],prg0[2556],prg0[2548],
                      prg0[2555],prg0[2547],prg0[2554],prg0[2546],prg0[2553],prg0[2545],prg0[2552],prg0[2544],
                      prg0[2543],prg0[2535],prg0[2542],prg0[2534],prg0[2541],prg0[2533],prg0[2540],prg0[2532],
                      prg0[2539],prg0[2531],prg0[2538],prg0[2530],prg0[2537],prg0[2529],prg0[2536],prg0[2528],
                      prg0[2527],prg0[2519],prg0[2526],prg0[2518],prg0[2525],prg0[2517],prg0[2524],prg0[2516],
                      prg0[2523],prg0[2515],prg0[2522],prg0[2514],prg0[2521],prg0[2513],prg0[2520],prg0[2512],
                      prg0[2511],prg0[2503],prg0[2510],prg0[2502],prg0[2509],prg0[2501],prg0[2508],prg0[2500],
                      prg0[2507],prg0[2499],prg0[2506],prg0[2498],prg0[2505],prg0[2497],prg0[2504],prg0[2496],
                      prg0[2495],prg0[2487],prg0[2494],prg0[2486],prg0[2493],prg0[2485],prg0[2492],prg0[2484],
                      prg0[2491],prg0[2483],prg0[2490],prg0[2482],prg0[2489],prg0[2481],prg0[2488],prg0[2480],
                      prg0[2479],prg0[2471],prg0[2478],prg0[2470],prg0[2477],prg0[2469],prg0[2476],prg0[2468],
                      prg0[2475],prg0[2467],prg0[2474],prg0[2466],prg0[2473],prg0[2465],prg0[2472],prg0[2464],
                      prg0[2463],prg0[2455],prg0[2462],prg0[2454],prg0[2461],prg0[2453],prg0[2460],prg0[2452],
                      prg0[2459],prg0[2451],prg0[2458],prg0[2450],prg0[2457],prg0[2449],prg0[2456],prg0[2448],
                      prg0[2447],prg0[2439],prg0[2446],prg0[2438],prg0[2445],prg0[2437],prg0[2444],prg0[2436],
                      prg0[2443],prg0[2435],prg0[2442],prg0[2434],prg0[2441],prg0[2433],prg0[2440],prg0[2432],
                      prg0[2431],prg0[2423],prg0[2430],prg0[2422],prg0[2429],prg0[2421],prg0[2428],prg0[2420],
                      prg0[2427],prg0[2419],prg0[2426],prg0[2418],prg0[2425],prg0[2417],prg0[2424],prg0[2416],
                      prg0[2415],prg0[2407],prg0[2414],prg0[2406],prg0[2413],prg0[2405],prg0[2412],prg0[2404],
                      prg0[2411],prg0[2403],prg0[2410],prg0[2402],prg0[2409],prg0[2401],prg0[2408],prg0[2400],
                      prg0[2399],prg0[2391],prg0[2398],prg0[2390],prg0[2397],prg0[2389],prg0[2396],prg0[2388],
                      prg0[2395],prg0[2387],prg0[2394],prg0[2386],prg0[2393],prg0[2385],prg0[2392],prg0[2384],
                      prg0[2383],prg0[2375],prg0[2382],prg0[2374],prg0[2381],prg0[2373],prg0[2380],prg0[2372],
                      prg0[2379],prg0[2371],prg0[2378],prg0[2370],prg0[2377],prg0[2369],prg0[2376],prg0[2368],
                      prg0[2367],prg0[2359],prg0[2366],prg0[2358],prg0[2365],prg0[2357],prg0[2364],prg0[2356],
                      prg0[2363],prg0[2355],prg0[2362],prg0[2354],prg0[2361],prg0[2353],prg0[2360],prg0[2352],
                      prg0[2351],prg0[2343],prg0[2350],prg0[2342],prg0[2349],prg0[2341],prg0[2348],prg0[2340],
                      prg0[2347],prg0[2339],prg0[2346],prg0[2338],prg0[2345],prg0[2337],prg0[2344],prg0[2336],
                      prg0[2335],prg0[2327],prg0[2334],prg0[2326],prg0[2333],prg0[2325],prg0[2332],prg0[2324],
                      prg0[2331],prg0[2323],prg0[2330],prg0[2322],prg0[2329],prg0[2321],prg0[2328],prg0[2320],
                      prg0[2319],prg0[2311],prg0[2318],prg0[2310],prg0[2317],prg0[2309],prg0[2316],prg0[2308],
                      prg0[2315],prg0[2307],prg0[2314],prg0[2306],prg0[2313],prg0[2305],prg0[2312],prg0[2304]}),
             .INIT_8({prg0[2303],prg0[2295],prg0[2302],prg0[2294],prg0[2301],prg0[2293],prg0[2300],prg0[2292],
                      prg0[2299],prg0[2291],prg0[2298],prg0[2290],prg0[2297],prg0[2289],prg0[2296],prg0[2288],
                      prg0[2287],prg0[2279],prg0[2286],prg0[2278],prg0[2285],prg0[2277],prg0[2284],prg0[2276],
                      prg0[2283],prg0[2275],prg0[2282],prg0[2274],prg0[2281],prg0[2273],prg0[2280],prg0[2272],
                      prg0[2271],prg0[2263],prg0[2270],prg0[2262],prg0[2269],prg0[2261],prg0[2268],prg0[2260],
                      prg0[2267],prg0[2259],prg0[2266],prg0[2258],prg0[2265],prg0[2257],prg0[2264],prg0[2256],
                      prg0[2255],prg0[2247],prg0[2254],prg0[2246],prg0[2253],prg0[2245],prg0[2252],prg0[2244],
                      prg0[2251],prg0[2243],prg0[2250],prg0[2242],prg0[2249],prg0[2241],prg0[2248],prg0[2240],
                      prg0[2239],prg0[2231],prg0[2238],prg0[2230],prg0[2237],prg0[2229],prg0[2236],prg0[2228],
                      prg0[2235],prg0[2227],prg0[2234],prg0[2226],prg0[2233],prg0[2225],prg0[2232],prg0[2224],
                      prg0[2223],prg0[2215],prg0[2222],prg0[2214],prg0[2221],prg0[2213],prg0[2220],prg0[2212],
                      prg0[2219],prg0[2211],prg0[2218],prg0[2210],prg0[2217],prg0[2209],prg0[2216],prg0[2208],
                      prg0[2207],prg0[2199],prg0[2206],prg0[2198],prg0[2205],prg0[2197],prg0[2204],prg0[2196],
                      prg0[2203],prg0[2195],prg0[2202],prg0[2194],prg0[2201],prg0[2193],prg0[2200],prg0[2192],
                      prg0[2191],prg0[2183],prg0[2190],prg0[2182],prg0[2189],prg0[2181],prg0[2188],prg0[2180],
                      prg0[2187],prg0[2179],prg0[2186],prg0[2178],prg0[2185],prg0[2177],prg0[2184],prg0[2176],
                      prg0[2175],prg0[2167],prg0[2174],prg0[2166],prg0[2173],prg0[2165],prg0[2172],prg0[2164],
                      prg0[2171],prg0[2163],prg0[2170],prg0[2162],prg0[2169],prg0[2161],prg0[2168],prg0[2160],
                      prg0[2159],prg0[2151],prg0[2158],prg0[2150],prg0[2157],prg0[2149],prg0[2156],prg0[2148],
                      prg0[2155],prg0[2147],prg0[2154],prg0[2146],prg0[2153],prg0[2145],prg0[2152],prg0[2144],
                      prg0[2143],prg0[2135],prg0[2142],prg0[2134],prg0[2141],prg0[2133],prg0[2140],prg0[2132],
                      prg0[2139],prg0[2131],prg0[2138],prg0[2130],prg0[2137],prg0[2129],prg0[2136],prg0[2128],
                      prg0[2127],prg0[2119],prg0[2126],prg0[2118],prg0[2125],prg0[2117],prg0[2124],prg0[2116],
                      prg0[2123],prg0[2115],prg0[2122],prg0[2114],prg0[2121],prg0[2113],prg0[2120],prg0[2112],
                      prg0[2111],prg0[2103],prg0[2110],prg0[2102],prg0[2109],prg0[2101],prg0[2108],prg0[2100],
                      prg0[2107],prg0[2099],prg0[2106],prg0[2098],prg0[2105],prg0[2097],prg0[2104],prg0[2096],
                      prg0[2095],prg0[2087],prg0[2094],prg0[2086],prg0[2093],prg0[2085],prg0[2092],prg0[2084],
                      prg0[2091],prg0[2083],prg0[2090],prg0[2082],prg0[2089],prg0[2081],prg0[2088],prg0[2080],
                      prg0[2079],prg0[2071],prg0[2078],prg0[2070],prg0[2077],prg0[2069],prg0[2076],prg0[2068],
                      prg0[2075],prg0[2067],prg0[2074],prg0[2066],prg0[2073],prg0[2065],prg0[2072],prg0[2064],
                      prg0[2063],prg0[2055],prg0[2062],prg0[2054],prg0[2061],prg0[2053],prg0[2060],prg0[2052],
                      prg0[2059],prg0[2051],prg0[2058],prg0[2050],prg0[2057],prg0[2049],prg0[2056],prg0[2048]}),
             .INIT_7({prg0[2047],prg0[2039],prg0[2046],prg0[2038],prg0[2045],prg0[2037],prg0[2044],prg0[2036],
                      prg0[2043],prg0[2035],prg0[2042],prg0[2034],prg0[2041],prg0[2033],prg0[2040],prg0[2032],
                      prg0[2031],prg0[2023],prg0[2030],prg0[2022],prg0[2029],prg0[2021],prg0[2028],prg0[2020],
                      prg0[2027],prg0[2019],prg0[2026],prg0[2018],prg0[2025],prg0[2017],prg0[2024],prg0[2016],
                      prg0[2015],prg0[2007],prg0[2014],prg0[2006],prg0[2013],prg0[2005],prg0[2012],prg0[2004],
                      prg0[2011],prg0[2003],prg0[2010],prg0[2002],prg0[2009],prg0[2001],prg0[2008],prg0[2000],
                      prg0[1999],prg0[1991],prg0[1998],prg0[1990],prg0[1997],prg0[1989],prg0[1996],prg0[1988],
                      prg0[1995],prg0[1987],prg0[1994],prg0[1986],prg0[1993],prg0[1985],prg0[1992],prg0[1984],
                      prg0[1983],prg0[1975],prg0[1982],prg0[1974],prg0[1981],prg0[1973],prg0[1980],prg0[1972],
                      prg0[1979],prg0[1971],prg0[1978],prg0[1970],prg0[1977],prg0[1969],prg0[1976],prg0[1968],
                      prg0[1967],prg0[1959],prg0[1966],prg0[1958],prg0[1965],prg0[1957],prg0[1964],prg0[1956],
                      prg0[1963],prg0[1955],prg0[1962],prg0[1954],prg0[1961],prg0[1953],prg0[1960],prg0[1952],
                      prg0[1951],prg0[1943],prg0[1950],prg0[1942],prg0[1949],prg0[1941],prg0[1948],prg0[1940],
                      prg0[1947],prg0[1939],prg0[1946],prg0[1938],prg0[1945],prg0[1937],prg0[1944],prg0[1936],
                      prg0[1935],prg0[1927],prg0[1934],prg0[1926],prg0[1933],prg0[1925],prg0[1932],prg0[1924],
                      prg0[1931],prg0[1923],prg0[1930],prg0[1922],prg0[1929],prg0[1921],prg0[1928],prg0[1920],
                      prg0[1919],prg0[1911],prg0[1918],prg0[1910],prg0[1917],prg0[1909],prg0[1916],prg0[1908],
                      prg0[1915],prg0[1907],prg0[1914],prg0[1906],prg0[1913],prg0[1905],prg0[1912],prg0[1904],
                      prg0[1903],prg0[1895],prg0[1902],prg0[1894],prg0[1901],prg0[1893],prg0[1900],prg0[1892],
                      prg0[1899],prg0[1891],prg0[1898],prg0[1890],prg0[1897],prg0[1889],prg0[1896],prg0[1888],
                      prg0[1887],prg0[1879],prg0[1886],prg0[1878],prg0[1885],prg0[1877],prg0[1884],prg0[1876],
                      prg0[1883],prg0[1875],prg0[1882],prg0[1874],prg0[1881],prg0[1873],prg0[1880],prg0[1872],
                      prg0[1871],prg0[1863],prg0[1870],prg0[1862],prg0[1869],prg0[1861],prg0[1868],prg0[1860],
                      prg0[1867],prg0[1859],prg0[1866],prg0[1858],prg0[1865],prg0[1857],prg0[1864],prg0[1856],
                      prg0[1855],prg0[1847],prg0[1854],prg0[1846],prg0[1853],prg0[1845],prg0[1852],prg0[1844],
                      prg0[1851],prg0[1843],prg0[1850],prg0[1842],prg0[1849],prg0[1841],prg0[1848],prg0[1840],
                      prg0[1839],prg0[1831],prg0[1838],prg0[1830],prg0[1837],prg0[1829],prg0[1836],prg0[1828],
                      prg0[1835],prg0[1827],prg0[1834],prg0[1826],prg0[1833],prg0[1825],prg0[1832],prg0[1824],
                      prg0[1823],prg0[1815],prg0[1822],prg0[1814],prg0[1821],prg0[1813],prg0[1820],prg0[1812],
                      prg0[1819],prg0[1811],prg0[1818],prg0[1810],prg0[1817],prg0[1809],prg0[1816],prg0[1808],
                      prg0[1807],prg0[1799],prg0[1806],prg0[1798],prg0[1805],prg0[1797],prg0[1804],prg0[1796],
                      prg0[1803],prg0[1795],prg0[1802],prg0[1794],prg0[1801],prg0[1793],prg0[1800],prg0[1792]}),
             .INIT_6({prg0[1791],prg0[1783],prg0[1790],prg0[1782],prg0[1789],prg0[1781],prg0[1788],prg0[1780],
                      prg0[1787],prg0[1779],prg0[1786],prg0[1778],prg0[1785],prg0[1777],prg0[1784],prg0[1776],
                      prg0[1775],prg0[1767],prg0[1774],prg0[1766],prg0[1773],prg0[1765],prg0[1772],prg0[1764],
                      prg0[1771],prg0[1763],prg0[1770],prg0[1762],prg0[1769],prg0[1761],prg0[1768],prg0[1760],
                      prg0[1759],prg0[1751],prg0[1758],prg0[1750],prg0[1757],prg0[1749],prg0[1756],prg0[1748],
                      prg0[1755],prg0[1747],prg0[1754],prg0[1746],prg0[1753],prg0[1745],prg0[1752],prg0[1744],
                      prg0[1743],prg0[1735],prg0[1742],prg0[1734],prg0[1741],prg0[1733],prg0[1740],prg0[1732],
                      prg0[1739],prg0[1731],prg0[1738],prg0[1730],prg0[1737],prg0[1729],prg0[1736],prg0[1728],
                      prg0[1727],prg0[1719],prg0[1726],prg0[1718],prg0[1725],prg0[1717],prg0[1724],prg0[1716],
                      prg0[1723],prg0[1715],prg0[1722],prg0[1714],prg0[1721],prg0[1713],prg0[1720],prg0[1712],
                      prg0[1711],prg0[1703],prg0[1710],prg0[1702],prg0[1709],prg0[1701],prg0[1708],prg0[1700],
                      prg0[1707],prg0[1699],prg0[1706],prg0[1698],prg0[1705],prg0[1697],prg0[1704],prg0[1696],
                      prg0[1695],prg0[1687],prg0[1694],prg0[1686],prg0[1693],prg0[1685],prg0[1692],prg0[1684],
                      prg0[1691],prg0[1683],prg0[1690],prg0[1682],prg0[1689],prg0[1681],prg0[1688],prg0[1680],
                      prg0[1679],prg0[1671],prg0[1678],prg0[1670],prg0[1677],prg0[1669],prg0[1676],prg0[1668],
                      prg0[1675],prg0[1667],prg0[1674],prg0[1666],prg0[1673],prg0[1665],prg0[1672],prg0[1664],
                      prg0[1663],prg0[1655],prg0[1662],prg0[1654],prg0[1661],prg0[1653],prg0[1660],prg0[1652],
                      prg0[1659],prg0[1651],prg0[1658],prg0[1650],prg0[1657],prg0[1649],prg0[1656],prg0[1648],
                      prg0[1647],prg0[1639],prg0[1646],prg0[1638],prg0[1645],prg0[1637],prg0[1644],prg0[1636],
                      prg0[1643],prg0[1635],prg0[1642],prg0[1634],prg0[1641],prg0[1633],prg0[1640],prg0[1632],
                      prg0[1631],prg0[1623],prg0[1630],prg0[1622],prg0[1629],prg0[1621],prg0[1628],prg0[1620],
                      prg0[1627],prg0[1619],prg0[1626],prg0[1618],prg0[1625],prg0[1617],prg0[1624],prg0[1616],
                      prg0[1615],prg0[1607],prg0[1614],prg0[1606],prg0[1613],prg0[1605],prg0[1612],prg0[1604],
                      prg0[1611],prg0[1603],prg0[1610],prg0[1602],prg0[1609],prg0[1601],prg0[1608],prg0[1600],
                      prg0[1599],prg0[1591],prg0[1598],prg0[1590],prg0[1597],prg0[1589],prg0[1596],prg0[1588],
                      prg0[1595],prg0[1587],prg0[1594],prg0[1586],prg0[1593],prg0[1585],prg0[1592],prg0[1584],
                      prg0[1583],prg0[1575],prg0[1582],prg0[1574],prg0[1581],prg0[1573],prg0[1580],prg0[1572],
                      prg0[1579],prg0[1571],prg0[1578],prg0[1570],prg0[1577],prg0[1569],prg0[1576],prg0[1568],
                      prg0[1567],prg0[1559],prg0[1566],prg0[1558],prg0[1565],prg0[1557],prg0[1564],prg0[1556],
                      prg0[1563],prg0[1555],prg0[1562],prg0[1554],prg0[1561],prg0[1553],prg0[1560],prg0[1552],
                      prg0[1551],prg0[1543],prg0[1550],prg0[1542],prg0[1549],prg0[1541],prg0[1548],prg0[1540],
                      prg0[1547],prg0[1539],prg0[1546],prg0[1538],prg0[1545],prg0[1537],prg0[1544],prg0[1536]}),
             .INIT_5({prg0[1535],prg0[1527],prg0[1534],prg0[1526],prg0[1533],prg0[1525],prg0[1532],prg0[1524],
                      prg0[1531],prg0[1523],prg0[1530],prg0[1522],prg0[1529],prg0[1521],prg0[1528],prg0[1520],
                      prg0[1519],prg0[1511],prg0[1518],prg0[1510],prg0[1517],prg0[1509],prg0[1516],prg0[1508],
                      prg0[1515],prg0[1507],prg0[1514],prg0[1506],prg0[1513],prg0[1505],prg0[1512],prg0[1504],
                      prg0[1503],prg0[1495],prg0[1502],prg0[1494],prg0[1501],prg0[1493],prg0[1500],prg0[1492],
                      prg0[1499],prg0[1491],prg0[1498],prg0[1490],prg0[1497],prg0[1489],prg0[1496],prg0[1488],
                      prg0[1487],prg0[1479],prg0[1486],prg0[1478],prg0[1485],prg0[1477],prg0[1484],prg0[1476],
                      prg0[1483],prg0[1475],prg0[1482],prg0[1474],prg0[1481],prg0[1473],prg0[1480],prg0[1472],
                      prg0[1471],prg0[1463],prg0[1470],prg0[1462],prg0[1469],prg0[1461],prg0[1468],prg0[1460],
                      prg0[1467],prg0[1459],prg0[1466],prg0[1458],prg0[1465],prg0[1457],prg0[1464],prg0[1456],
                      prg0[1455],prg0[1447],prg0[1454],prg0[1446],prg0[1453],prg0[1445],prg0[1452],prg0[1444],
                      prg0[1451],prg0[1443],prg0[1450],prg0[1442],prg0[1449],prg0[1441],prg0[1448],prg0[1440],
                      prg0[1439],prg0[1431],prg0[1438],prg0[1430],prg0[1437],prg0[1429],prg0[1436],prg0[1428],
                      prg0[1435],prg0[1427],prg0[1434],prg0[1426],prg0[1433],prg0[1425],prg0[1432],prg0[1424],
                      prg0[1423],prg0[1415],prg0[1422],prg0[1414],prg0[1421],prg0[1413],prg0[1420],prg0[1412],
                      prg0[1419],prg0[1411],prg0[1418],prg0[1410],prg0[1417],prg0[1409],prg0[1416],prg0[1408],
                      prg0[1407],prg0[1399],prg0[1406],prg0[1398],prg0[1405],prg0[1397],prg0[1404],prg0[1396],
                      prg0[1403],prg0[1395],prg0[1402],prg0[1394],prg0[1401],prg0[1393],prg0[1400],prg0[1392],
                      prg0[1391],prg0[1383],prg0[1390],prg0[1382],prg0[1389],prg0[1381],prg0[1388],prg0[1380],
                      prg0[1387],prg0[1379],prg0[1386],prg0[1378],prg0[1385],prg0[1377],prg0[1384],prg0[1376],
                      prg0[1375],prg0[1367],prg0[1374],prg0[1366],prg0[1373],prg0[1365],prg0[1372],prg0[1364],
                      prg0[1371],prg0[1363],prg0[1370],prg0[1362],prg0[1369],prg0[1361],prg0[1368],prg0[1360],
                      prg0[1359],prg0[1351],prg0[1358],prg0[1350],prg0[1357],prg0[1349],prg0[1356],prg0[1348],
                      prg0[1355],prg0[1347],prg0[1354],prg0[1346],prg0[1353],prg0[1345],prg0[1352],prg0[1344],
                      prg0[1343],prg0[1335],prg0[1342],prg0[1334],prg0[1341],prg0[1333],prg0[1340],prg0[1332],
                      prg0[1339],prg0[1331],prg0[1338],prg0[1330],prg0[1337],prg0[1329],prg0[1336],prg0[1328],
                      prg0[1327],prg0[1319],prg0[1326],prg0[1318],prg0[1325],prg0[1317],prg0[1324],prg0[1316],
                      prg0[1323],prg0[1315],prg0[1322],prg0[1314],prg0[1321],prg0[1313],prg0[1320],prg0[1312],
                      prg0[1311],prg0[1303],prg0[1310],prg0[1302],prg0[1309],prg0[1301],prg0[1308],prg0[1300],
                      prg0[1307],prg0[1299],prg0[1306],prg0[1298],prg0[1305],prg0[1297],prg0[1304],prg0[1296],
                      prg0[1295],prg0[1287],prg0[1294],prg0[1286],prg0[1293],prg0[1285],prg0[1292],prg0[1284],
                      prg0[1291],prg0[1283],prg0[1290],prg0[1282],prg0[1289],prg0[1281],prg0[1288],prg0[1280]}),
             .INIT_4({prg0[1279],prg0[1271],prg0[1278],prg0[1270],prg0[1277],prg0[1269],prg0[1276],prg0[1268],
                      prg0[1275],prg0[1267],prg0[1274],prg0[1266],prg0[1273],prg0[1265],prg0[1272],prg0[1264],
                      prg0[1263],prg0[1255],prg0[1262],prg0[1254],prg0[1261],prg0[1253],prg0[1260],prg0[1252],
                      prg0[1259],prg0[1251],prg0[1258],prg0[1250],prg0[1257],prg0[1249],prg0[1256],prg0[1248],
                      prg0[1247],prg0[1239],prg0[1246],prg0[1238],prg0[1245],prg0[1237],prg0[1244],prg0[1236],
                      prg0[1243],prg0[1235],prg0[1242],prg0[1234],prg0[1241],prg0[1233],prg0[1240],prg0[1232],
                      prg0[1231],prg0[1223],prg0[1230],prg0[1222],prg0[1229],prg0[1221],prg0[1228],prg0[1220],
                      prg0[1227],prg0[1219],prg0[1226],prg0[1218],prg0[1225],prg0[1217],prg0[1224],prg0[1216],
                      prg0[1215],prg0[1207],prg0[1214],prg0[1206],prg0[1213],prg0[1205],prg0[1212],prg0[1204],
                      prg0[1211],prg0[1203],prg0[1210],prg0[1202],prg0[1209],prg0[1201],prg0[1208],prg0[1200],
                      prg0[1199],prg0[1191],prg0[1198],prg0[1190],prg0[1197],prg0[1189],prg0[1196],prg0[1188],
                      prg0[1195],prg0[1187],prg0[1194],prg0[1186],prg0[1193],prg0[1185],prg0[1192],prg0[1184],
                      prg0[1183],prg0[1175],prg0[1182],prg0[1174],prg0[1181],prg0[1173],prg0[1180],prg0[1172],
                      prg0[1179],prg0[1171],prg0[1178],prg0[1170],prg0[1177],prg0[1169],prg0[1176],prg0[1168],
                      prg0[1167],prg0[1159],prg0[1166],prg0[1158],prg0[1165],prg0[1157],prg0[1164],prg0[1156],
                      prg0[1163],prg0[1155],prg0[1162],prg0[1154],prg0[1161],prg0[1153],prg0[1160],prg0[1152],
                      prg0[1151],prg0[1143],prg0[1150],prg0[1142],prg0[1149],prg0[1141],prg0[1148],prg0[1140],
                      prg0[1147],prg0[1139],prg0[1146],prg0[1138],prg0[1145],prg0[1137],prg0[1144],prg0[1136],
                      prg0[1135],prg0[1127],prg0[1134],prg0[1126],prg0[1133],prg0[1125],prg0[1132],prg0[1124],
                      prg0[1131],prg0[1123],prg0[1130],prg0[1122],prg0[1129],prg0[1121],prg0[1128],prg0[1120],
                      prg0[1119],prg0[1111],prg0[1118],prg0[1110],prg0[1117],prg0[1109],prg0[1116],prg0[1108],
                      prg0[1115],prg0[1107],prg0[1114],prg0[1106],prg0[1113],prg0[1105],prg0[1112],prg0[1104],
                      prg0[1103],prg0[1095],prg0[1102],prg0[1094],prg0[1101],prg0[1093],prg0[1100],prg0[1092],
                      prg0[1099],prg0[1091],prg0[1098],prg0[1090],prg0[1097],prg0[1089],prg0[1096],prg0[1088],
                      prg0[1087],prg0[1079],prg0[1086],prg0[1078],prg0[1085],prg0[1077],prg0[1084],prg0[1076],
                      prg0[1083],prg0[1075],prg0[1082],prg0[1074],prg0[1081],prg0[1073],prg0[1080],prg0[1072],
                      prg0[1071],prg0[1063],prg0[1070],prg0[1062],prg0[1069],prg0[1061],prg0[1068],prg0[1060],
                      prg0[1067],prg0[1059],prg0[1066],prg0[1058],prg0[1065],prg0[1057],prg0[1064],prg0[1056],
                      prg0[1055],prg0[1047],prg0[1054],prg0[1046],prg0[1053],prg0[1045],prg0[1052],prg0[1044],
                      prg0[1051],prg0[1043],prg0[1050],prg0[1042],prg0[1049],prg0[1041],prg0[1048],prg0[1040],
                      prg0[1039],prg0[1031],prg0[1038],prg0[1030],prg0[1037],prg0[1029],prg0[1036],prg0[1028],
                      prg0[1035],prg0[1027],prg0[1034],prg0[1026],prg0[1033],prg0[1025],prg0[1032],prg0[1024]}),
             .INIT_3({prg0[1023],prg0[1015],prg0[1022],prg0[1014],prg0[1021],prg0[1013],prg0[1020],prg0[1012],
                      prg0[1019],prg0[1011],prg0[1018],prg0[1010],prg0[1017],prg0[1009],prg0[1016],prg0[1008],
                      prg0[1007],prg0[ 999],prg0[1006],prg0[ 998],prg0[1005],prg0[ 997],prg0[1004],prg0[ 996],
                      prg0[1003],prg0[ 995],prg0[1002],prg0[ 994],prg0[1001],prg0[ 993],prg0[1000],prg0[ 992],
                      prg0[ 991],prg0[ 983],prg0[ 990],prg0[ 982],prg0[ 989],prg0[ 981],prg0[ 988],prg0[ 980],
                      prg0[ 987],prg0[ 979],prg0[ 986],prg0[ 978],prg0[ 985],prg0[ 977],prg0[ 984],prg0[ 976],
                      prg0[ 975],prg0[ 967],prg0[ 974],prg0[ 966],prg0[ 973],prg0[ 965],prg0[ 972],prg0[ 964],
                      prg0[ 971],prg0[ 963],prg0[ 970],prg0[ 962],prg0[ 969],prg0[ 961],prg0[ 968],prg0[ 960],
                      prg0[ 959],prg0[ 951],prg0[ 958],prg0[ 950],prg0[ 957],prg0[ 949],prg0[ 956],prg0[ 948],
                      prg0[ 955],prg0[ 947],prg0[ 954],prg0[ 946],prg0[ 953],prg0[ 945],prg0[ 952],prg0[ 944],
                      prg0[ 943],prg0[ 935],prg0[ 942],prg0[ 934],prg0[ 941],prg0[ 933],prg0[ 940],prg0[ 932],
                      prg0[ 939],prg0[ 931],prg0[ 938],prg0[ 930],prg0[ 937],prg0[ 929],prg0[ 936],prg0[ 928],
                      prg0[ 927],prg0[ 919],prg0[ 926],prg0[ 918],prg0[ 925],prg0[ 917],prg0[ 924],prg0[ 916],
                      prg0[ 923],prg0[ 915],prg0[ 922],prg0[ 914],prg0[ 921],prg0[ 913],prg0[ 920],prg0[ 912],
                      prg0[ 911],prg0[ 903],prg0[ 910],prg0[ 902],prg0[ 909],prg0[ 901],prg0[ 908],prg0[ 900],
                      prg0[ 907],prg0[ 899],prg0[ 906],prg0[ 898],prg0[ 905],prg0[ 897],prg0[ 904],prg0[ 896],
                      prg0[ 895],prg0[ 887],prg0[ 894],prg0[ 886],prg0[ 893],prg0[ 885],prg0[ 892],prg0[ 884],
                      prg0[ 891],prg0[ 883],prg0[ 890],prg0[ 882],prg0[ 889],prg0[ 881],prg0[ 888],prg0[ 880],
                      prg0[ 879],prg0[ 871],prg0[ 878],prg0[ 870],prg0[ 877],prg0[ 869],prg0[ 876],prg0[ 868],
                      prg0[ 875],prg0[ 867],prg0[ 874],prg0[ 866],prg0[ 873],prg0[ 865],prg0[ 872],prg0[ 864],
                      prg0[ 863],prg0[ 855],prg0[ 862],prg0[ 854],prg0[ 861],prg0[ 853],prg0[ 860],prg0[ 852],
                      prg0[ 859],prg0[ 851],prg0[ 858],prg0[ 850],prg0[ 857],prg0[ 849],prg0[ 856],prg0[ 848],
                      prg0[ 847],prg0[ 839],prg0[ 846],prg0[ 838],prg0[ 845],prg0[ 837],prg0[ 844],prg0[ 836],
                      prg0[ 843],prg0[ 835],prg0[ 842],prg0[ 834],prg0[ 841],prg0[ 833],prg0[ 840],prg0[ 832],
                      prg0[ 831],prg0[ 823],prg0[ 830],prg0[ 822],prg0[ 829],prg0[ 821],prg0[ 828],prg0[ 820],
                      prg0[ 827],prg0[ 819],prg0[ 826],prg0[ 818],prg0[ 825],prg0[ 817],prg0[ 824],prg0[ 816],
                      prg0[ 815],prg0[ 807],prg0[ 814],prg0[ 806],prg0[ 813],prg0[ 805],prg0[ 812],prg0[ 804],
                      prg0[ 811],prg0[ 803],prg0[ 810],prg0[ 802],prg0[ 809],prg0[ 801],prg0[ 808],prg0[ 800],
                      prg0[ 799],prg0[ 791],prg0[ 798],prg0[ 790],prg0[ 797],prg0[ 789],prg0[ 796],prg0[ 788],
                      prg0[ 795],prg0[ 787],prg0[ 794],prg0[ 786],prg0[ 793],prg0[ 785],prg0[ 792],prg0[ 784],
                      prg0[ 783],prg0[ 775],prg0[ 782],prg0[ 774],prg0[ 781],prg0[ 773],prg0[ 780],prg0[ 772],
                      prg0[ 779],prg0[ 771],prg0[ 778],prg0[ 770],prg0[ 777],prg0[ 769],prg0[ 776],prg0[ 768]}),
             .INIT_2({prg0[ 767],prg0[ 759],prg0[ 766],prg0[ 758],prg0[ 765],prg0[ 757],prg0[ 764],prg0[ 756],
                      prg0[ 763],prg0[ 755],prg0[ 762],prg0[ 754],prg0[ 761],prg0[ 753],prg0[ 760],prg0[ 752],
                      prg0[ 751],prg0[ 743],prg0[ 750],prg0[ 742],prg0[ 749],prg0[ 741],prg0[ 748],prg0[ 740],
                      prg0[ 747],prg0[ 739],prg0[ 746],prg0[ 738],prg0[ 745],prg0[ 737],prg0[ 744],prg0[ 736],
                      prg0[ 735],prg0[ 727],prg0[ 734],prg0[ 726],prg0[ 733],prg0[ 725],prg0[ 732],prg0[ 724],
                      prg0[ 731],prg0[ 723],prg0[ 730],prg0[ 722],prg0[ 729],prg0[ 721],prg0[ 728],prg0[ 720],
                      prg0[ 719],prg0[ 711],prg0[ 718],prg0[ 710],prg0[ 717],prg0[ 709],prg0[ 716],prg0[ 708],
                      prg0[ 715],prg0[ 707],prg0[ 714],prg0[ 706],prg0[ 713],prg0[ 705],prg0[ 712],prg0[ 704],
                      prg0[ 703],prg0[ 695],prg0[ 702],prg0[ 694],prg0[ 701],prg0[ 693],prg0[ 700],prg0[ 692],
                      prg0[ 699],prg0[ 691],prg0[ 698],prg0[ 690],prg0[ 697],prg0[ 689],prg0[ 696],prg0[ 688],
                      prg0[ 687],prg0[ 679],prg0[ 686],prg0[ 678],prg0[ 685],prg0[ 677],prg0[ 684],prg0[ 676],
                      prg0[ 683],prg0[ 675],prg0[ 682],prg0[ 674],prg0[ 681],prg0[ 673],prg0[ 680],prg0[ 672],
                      prg0[ 671],prg0[ 663],prg0[ 670],prg0[ 662],prg0[ 669],prg0[ 661],prg0[ 668],prg0[ 660],
                      prg0[ 667],prg0[ 659],prg0[ 666],prg0[ 658],prg0[ 665],prg0[ 657],prg0[ 664],prg0[ 656],
                      prg0[ 655],prg0[ 647],prg0[ 654],prg0[ 646],prg0[ 653],prg0[ 645],prg0[ 652],prg0[ 644],
                      prg0[ 651],prg0[ 643],prg0[ 650],prg0[ 642],prg0[ 649],prg0[ 641],prg0[ 648],prg0[ 640],
                      prg0[ 639],prg0[ 631],prg0[ 638],prg0[ 630],prg0[ 637],prg0[ 629],prg0[ 636],prg0[ 628],
                      prg0[ 635],prg0[ 627],prg0[ 634],prg0[ 626],prg0[ 633],prg0[ 625],prg0[ 632],prg0[ 624],
                      prg0[ 623],prg0[ 615],prg0[ 622],prg0[ 614],prg0[ 621],prg0[ 613],prg0[ 620],prg0[ 612],
                      prg0[ 619],prg0[ 611],prg0[ 618],prg0[ 610],prg0[ 617],prg0[ 609],prg0[ 616],prg0[ 608],
                      prg0[ 607],prg0[ 599],prg0[ 606],prg0[ 598],prg0[ 605],prg0[ 597],prg0[ 604],prg0[ 596],
                      prg0[ 603],prg0[ 595],prg0[ 602],prg0[ 594],prg0[ 601],prg0[ 593],prg0[ 600],prg0[ 592],
                      prg0[ 591],prg0[ 583],prg0[ 590],prg0[ 582],prg0[ 589],prg0[ 581],prg0[ 588],prg0[ 580],
                      prg0[ 587],prg0[ 579],prg0[ 586],prg0[ 578],prg0[ 585],prg0[ 577],prg0[ 584],prg0[ 576],
                      prg0[ 575],prg0[ 567],prg0[ 574],prg0[ 566],prg0[ 573],prg0[ 565],prg0[ 572],prg0[ 564],
                      prg0[ 571],prg0[ 563],prg0[ 570],prg0[ 562],prg0[ 569],prg0[ 561],prg0[ 568],prg0[ 560],
                      prg0[ 559],prg0[ 551],prg0[ 558],prg0[ 550],prg0[ 557],prg0[ 549],prg0[ 556],prg0[ 548],
                      prg0[ 555],prg0[ 547],prg0[ 554],prg0[ 546],prg0[ 553],prg0[ 545],prg0[ 552],prg0[ 544],
                      prg0[ 543],prg0[ 535],prg0[ 542],prg0[ 534],prg0[ 541],prg0[ 533],prg0[ 540],prg0[ 532],
                      prg0[ 539],prg0[ 531],prg0[ 538],prg0[ 530],prg0[ 537],prg0[ 529],prg0[ 536],prg0[ 528],
                      prg0[ 527],prg0[ 519],prg0[ 526],prg0[ 518],prg0[ 525],prg0[ 517],prg0[ 524],prg0[ 516],
                      prg0[ 523],prg0[ 515],prg0[ 522],prg0[ 514],prg0[ 521],prg0[ 513],prg0[ 520],prg0[ 512]}),
             .INIT_1({prg0[ 511],prg0[ 503],prg0[ 510],prg0[ 502],prg0[ 509],prg0[ 501],prg0[ 508],prg0[ 500],
                      prg0[ 507],prg0[ 499],prg0[ 506],prg0[ 498],prg0[ 505],prg0[ 497],prg0[ 504],prg0[ 496],
                      prg0[ 495],prg0[ 487],prg0[ 494],prg0[ 486],prg0[ 493],prg0[ 485],prg0[ 492],prg0[ 484],
                      prg0[ 491],prg0[ 483],prg0[ 490],prg0[ 482],prg0[ 489],prg0[ 481],prg0[ 488],prg0[ 480],
                      prg0[ 479],prg0[ 471],prg0[ 478],prg0[ 470],prg0[ 477],prg0[ 469],prg0[ 476],prg0[ 468],
                      prg0[ 475],prg0[ 467],prg0[ 474],prg0[ 466],prg0[ 473],prg0[ 465],prg0[ 472],prg0[ 464],
                      prg0[ 463],prg0[ 455],prg0[ 462],prg0[ 454],prg0[ 461],prg0[ 453],prg0[ 460],prg0[ 452],
                      prg0[ 459],prg0[ 451],prg0[ 458],prg0[ 450],prg0[ 457],prg0[ 449],prg0[ 456],prg0[ 448],
                      prg0[ 447],prg0[ 439],prg0[ 446],prg0[ 438],prg0[ 445],prg0[ 437],prg0[ 444],prg0[ 436],
                      prg0[ 443],prg0[ 435],prg0[ 442],prg0[ 434],prg0[ 441],prg0[ 433],prg0[ 440],prg0[ 432],
                      prg0[ 431],prg0[ 423],prg0[ 430],prg0[ 422],prg0[ 429],prg0[ 421],prg0[ 428],prg0[ 420],
                      prg0[ 427],prg0[ 419],prg0[ 426],prg0[ 418],prg0[ 425],prg0[ 417],prg0[ 424],prg0[ 416],
                      prg0[ 415],prg0[ 407],prg0[ 414],prg0[ 406],prg0[ 413],prg0[ 405],prg0[ 412],prg0[ 404],
                      prg0[ 411],prg0[ 403],prg0[ 410],prg0[ 402],prg0[ 409],prg0[ 401],prg0[ 408],prg0[ 400],
                      prg0[ 399],prg0[ 391],prg0[ 398],prg0[ 390],prg0[ 397],prg0[ 389],prg0[ 396],prg0[ 388],
                      prg0[ 395],prg0[ 387],prg0[ 394],prg0[ 386],prg0[ 393],prg0[ 385],prg0[ 392],prg0[ 384],
                      prg0[ 383],prg0[ 375],prg0[ 382],prg0[ 374],prg0[ 381],prg0[ 373],prg0[ 380],prg0[ 372],
                      prg0[ 379],prg0[ 371],prg0[ 378],prg0[ 370],prg0[ 377],prg0[ 369],prg0[ 376],prg0[ 368],
                      prg0[ 367],prg0[ 359],prg0[ 366],prg0[ 358],prg0[ 365],prg0[ 357],prg0[ 364],prg0[ 356],
                      prg0[ 363],prg0[ 355],prg0[ 362],prg0[ 354],prg0[ 361],prg0[ 353],prg0[ 360],prg0[ 352],
                      prg0[ 351],prg0[ 343],prg0[ 350],prg0[ 342],prg0[ 349],prg0[ 341],prg0[ 348],prg0[ 340],
                      prg0[ 347],prg0[ 339],prg0[ 346],prg0[ 338],prg0[ 345],prg0[ 337],prg0[ 344],prg0[ 336],
                      prg0[ 335],prg0[ 327],prg0[ 334],prg0[ 326],prg0[ 333],prg0[ 325],prg0[ 332],prg0[ 324],
                      prg0[ 331],prg0[ 323],prg0[ 330],prg0[ 322],prg0[ 329],prg0[ 321],prg0[ 328],prg0[ 320],
                      prg0[ 319],prg0[ 311],prg0[ 318],prg0[ 310],prg0[ 317],prg0[ 309],prg0[ 316],prg0[ 308],
                      prg0[ 315],prg0[ 307],prg0[ 314],prg0[ 306],prg0[ 313],prg0[ 305],prg0[ 312],prg0[ 304],
                      prg0[ 303],prg0[ 295],prg0[ 302],prg0[ 294],prg0[ 301],prg0[ 293],prg0[ 300],prg0[ 292],
                      prg0[ 299],prg0[ 291],prg0[ 298],prg0[ 290],prg0[ 297],prg0[ 289],prg0[ 296],prg0[ 288],
                      prg0[ 287],prg0[ 279],prg0[ 286],prg0[ 278],prg0[ 285],prg0[ 277],prg0[ 284],prg0[ 276],
                      prg0[ 283],prg0[ 275],prg0[ 282],prg0[ 274],prg0[ 281],prg0[ 273],prg0[ 280],prg0[ 272],
                      prg0[ 271],prg0[ 263],prg0[ 270],prg0[ 262],prg0[ 269],prg0[ 261],prg0[ 268],prg0[ 260],
                      prg0[ 267],prg0[ 259],prg0[ 266],prg0[ 258],prg0[ 265],prg0[ 257],prg0[ 264],prg0[ 256]}),
             .INIT_0({prg0[ 255],prg0[ 247],prg0[ 254],prg0[ 246],prg0[ 253],prg0[ 245],prg0[ 252],prg0[ 244],
                      prg0[ 251],prg0[ 243],prg0[ 250],prg0[ 242],prg0[ 249],prg0[ 241],prg0[ 248],prg0[ 240],
                      prg0[ 239],prg0[ 231],prg0[ 238],prg0[ 230],prg0[ 237],prg0[ 229],prg0[ 236],prg0[ 228],
                      prg0[ 235],prg0[ 227],prg0[ 234],prg0[ 226],prg0[ 233],prg0[ 225],prg0[ 232],prg0[ 224],
                      prg0[ 223],prg0[ 215],prg0[ 222],prg0[ 214],prg0[ 221],prg0[ 213],prg0[ 220],prg0[ 212],
                      prg0[ 219],prg0[ 211],prg0[ 218],prg0[ 210],prg0[ 217],prg0[ 209],prg0[ 216],prg0[ 208],
                      prg0[ 207],prg0[ 199],prg0[ 206],prg0[ 198],prg0[ 205],prg0[ 197],prg0[ 204],prg0[ 196],
                      prg0[ 203],prg0[ 195],prg0[ 202],prg0[ 194],prg0[ 201],prg0[ 193],prg0[ 200],prg0[ 192],
                      prg0[ 191],prg0[ 183],prg0[ 190],prg0[ 182],prg0[ 189],prg0[ 181],prg0[ 188],prg0[ 180],
                      prg0[ 187],prg0[ 179],prg0[ 186],prg0[ 178],prg0[ 185],prg0[ 177],prg0[ 184],prg0[ 176],
                      prg0[ 175],prg0[ 167],prg0[ 174],prg0[ 166],prg0[ 173],prg0[ 165],prg0[ 172],prg0[ 164],
                      prg0[ 171],prg0[ 163],prg0[ 170],prg0[ 162],prg0[ 169],prg0[ 161],prg0[ 168],prg0[ 160],
                      prg0[ 159],prg0[ 151],prg0[ 158],prg0[ 150],prg0[ 157],prg0[ 149],prg0[ 156],prg0[ 148],
                      prg0[ 155],prg0[ 147],prg0[ 154],prg0[ 146],prg0[ 153],prg0[ 145],prg0[ 152],prg0[ 144],
                      prg0[ 143],prg0[ 135],prg0[ 142],prg0[ 134],prg0[ 141],prg0[ 133],prg0[ 140],prg0[ 132],
                      prg0[ 139],prg0[ 131],prg0[ 138],prg0[ 130],prg0[ 137],prg0[ 129],prg0[ 136],prg0[ 128],
                      prg0[ 127],prg0[ 119],prg0[ 126],prg0[ 118],prg0[ 125],prg0[ 117],prg0[ 124],prg0[ 116],
                      prg0[ 123],prg0[ 115],prg0[ 122],prg0[ 114],prg0[ 121],prg0[ 113],prg0[ 120],prg0[ 112],
                      prg0[ 111],prg0[ 103],prg0[ 110],prg0[ 102],prg0[ 109],prg0[ 101],prg0[ 108],prg0[ 100],
                      prg0[ 107],prg0[  99],prg0[ 106],prg0[  98],prg0[ 105],prg0[  97],prg0[ 104],prg0[  96],
                      prg0[  95],prg0[  87],prg0[  94],prg0[  86],prg0[  93],prg0[  85],prg0[  92],prg0[  84],
                      prg0[  91],prg0[  83],prg0[  90],prg0[  82],prg0[  89],prg0[  81],prg0[  88],prg0[  80],
                      prg0[  79],prg0[  71],prg0[  78],prg0[  70],prg0[  77],prg0[  69],prg0[  76],prg0[  68],
                      prg0[  75],prg0[  67],prg0[  74],prg0[  66],prg0[  73],prg0[  65],prg0[  72],prg0[  64],
                      prg0[  63],prg0[  55],prg0[  62],prg0[  54],prg0[  61],prg0[  53],prg0[  60],prg0[  52],
                      prg0[  59],prg0[  51],prg0[  58],prg0[  50],prg0[  57],prg0[  49],prg0[  56],prg0[  48],
                      prg0[  47],prg0[  39],prg0[  46],prg0[  38],prg0[  45],prg0[  37],prg0[  44],prg0[  36],
                      prg0[  43],prg0[  35],prg0[  42],prg0[  34],prg0[  41],prg0[  33],prg0[  40],prg0[  32],
                      prg0[  31],prg0[  23],prg0[  30],prg0[  22],prg0[  29],prg0[  21],prg0[  28],prg0[  20],
                      prg0[  27],prg0[  19],prg0[  26],prg0[  18],prg0[  25],prg0[  17],prg0[  24],prg0[  16],
                      prg0[  15],prg0[   7],prg0[  14],prg0[   6],prg0[  13],prg0[   5],prg0[  12],prg0[   4],
                      prg0[  11],prg0[   3],prg0[  10],prg0[   2],prg0[   9],prg0[   1],prg0[   8],prg0[   0]}),
             .READ_MODE(1),
             .WRITE_MODE(1))
         mem
           (// Outputs
            .RDATA  ( {dum8[7],DAT_O[7],
                       dum8[6],DAT_O[6],
                       dum8[5],DAT_O[5],
                       dum8[4],DAT_O[4],
                       dum8[3],DAT_O[3],
                       dum8[2],DAT_O[2],
                       dum8[1],DAT_O[1],
                       dum8[0],DAT_O[0]}            ),
            // Input
            .MASK   ( 16'h0                         ),
            .WDATA  ( {1'b0, B[7],1'b0, B[6],
                       1'b0, B[5],1'b0, B[4],
                       1'b0, B[3],1'b0, B[2],
                       1'b0, B[1],1'b0, B[0]}       ),                       
            .WADDR  ( {2'b0,Wai[0],Wai[8:1]}        ), // Note mangling
            .RADDR  ( {2'b0,Rai[0],Rai[8:1]}        ), // Note mangling
            .RE     ( 1'b1                          ),
            .WE     ( we                            ), // May perhaps save a lut. use .WE(iwe) .WCLKE(~bmask)
            .WCLK   ( clk                           ),
            .RCLK   ( clk                           ),
            .RCLKE  ( 1'b1                          ),
            .WCLKE  ( 1'b1                          ) //  May perhaps save a lut. use .WE(iwe) .WCLKE(~bmask)
            /*AUTOINST*/);
         
      end else begin
         /* Split up to 2 KiB memory into low and high nibbles
          */
         localparam [4095:0]
           pb1 = {prg3[4091:4088],prg3[4083:4080],prg3[4075:4072],prg3[4067:4064],prg3[4059:4056],prg3[4051:4048],prg3[4043:4040],prg3[4035:4032],
                  prg3[4027:4024],prg3[4019:4016],prg3[4011:4008],prg3[4003:4000],prg3[3995:3992],prg3[3987:3984],prg3[3979:3976],prg3[3971:3968],
                  prg3[3963:3960],prg3[3955:3952],prg3[3947:3944],prg3[3939:3936],prg3[3931:3928],prg3[3923:3920],prg3[3915:3912],prg3[3907:3904],
                  prg3[3899:3896],prg3[3891:3888],prg3[3883:3880],prg3[3875:3872],prg3[3867:3864],prg3[3859:3856],prg3[3851:3848],prg3[3843:3840],
                  prg3[3835:3832],prg3[3827:3824],prg3[3819:3816],prg3[3811:3808],prg3[3803:3800],prg3[3795:3792],prg3[3787:3784],prg3[3779:3776],
                  prg3[3771:3768],prg3[3763:3760],prg3[3755:3752],prg3[3747:3744],prg3[3739:3736],prg3[3731:3728],prg3[3723:3720],prg3[3715:3712],
                  prg3[3707:3704],prg3[3699:3696],prg3[3691:3688],prg3[3683:3680],prg3[3675:3672],prg3[3667:3664],prg3[3659:3656],prg3[3651:3648],
                  prg3[3643:3640],prg3[3635:3632],prg3[3627:3624],prg3[3619:3616],prg3[3611:3608],prg3[3603:3600],prg3[3595:3592],prg3[3587:3584],
                  prg3[3579:3576],prg3[3571:3568],prg3[3563:3560],prg3[3555:3552],prg3[3547:3544],prg3[3539:3536],prg3[3531:3528],prg3[3523:3520],
                  prg3[3515:3512],prg3[3507:3504],prg3[3499:3496],prg3[3491:3488],prg3[3483:3480],prg3[3475:3472],prg3[3467:3464],prg3[3459:3456],
                  prg3[3451:3448],prg3[3443:3440],prg3[3435:3432],prg3[3427:3424],prg3[3419:3416],prg3[3411:3408],prg3[3403:3400],prg3[3395:3392],
                  prg3[3387:3384],prg3[3379:3376],prg3[3371:3368],prg3[3363:3360],prg3[3355:3352],prg3[3347:3344],prg3[3339:3336],prg3[3331:3328],
                  prg3[3323:3320],prg3[3315:3312],prg3[3307:3304],prg3[3299:3296],prg3[3291:3288],prg3[3283:3280],prg3[3275:3272],prg3[3267:3264],
                  prg3[3259:3256],prg3[3251:3248],prg3[3243:3240],prg3[3235:3232],prg3[3227:3224],prg3[3219:3216],prg3[3211:3208],prg3[3203:3200],
                  prg3[3195:3192],prg3[3187:3184],prg3[3179:3176],prg3[3171:3168],prg3[3163:3160],prg3[3155:3152],prg3[3147:3144],prg3[3139:3136],
                  prg3[3131:3128],prg3[3123:3120],prg3[3115:3112],prg3[3107:3104],prg3[3099:3096],prg3[3091:3088],prg3[3083:3080],prg3[3075:3072],
                  prg3[3067:3064],prg3[3059:3056],prg3[3051:3048],prg3[3043:3040],prg3[3035:3032],prg3[3027:3024],prg3[3019:3016],prg3[3011:3008],
                  prg3[3003:3000],prg3[2995:2992],prg3[2987:2984],prg3[2979:2976],prg3[2971:2968],prg3[2963:2960],prg3[2955:2952],prg3[2947:2944],
                  prg3[2939:2936],prg3[2931:2928],prg3[2923:2920],prg3[2915:2912],prg3[2907:2904],prg3[2899:2896],prg3[2891:2888],prg3[2883:2880],
                  prg3[2875:2872],prg3[2867:2864],prg3[2859:2856],prg3[2851:2848],prg3[2843:2840],prg3[2835:2832],prg3[2827:2824],prg3[2819:2816],
                  prg3[2811:2808],prg3[2803:2800],prg3[2795:2792],prg3[2787:2784],prg3[2779:2776],prg3[2771:2768],prg3[2763:2760],prg3[2755:2752],
                  prg3[2747:2744],prg3[2739:2736],prg3[2731:2728],prg3[2723:2720],prg3[2715:2712],prg3[2707:2704],prg3[2699:2696],prg3[2691:2688],
                  prg3[2683:2680],prg3[2675:2672],prg3[2667:2664],prg3[2659:2656],prg3[2651:2648],prg3[2643:2640],prg3[2635:2632],prg3[2627:2624],
                  prg3[2619:2616],prg3[2611:2608],prg3[2603:2600],prg3[2595:2592],prg3[2587:2584],prg3[2579:2576],prg3[2571:2568],prg3[2563:2560],
                  prg3[2555:2552],prg3[2547:2544],prg3[2539:2536],prg3[2531:2528],prg3[2523:2520],prg3[2515:2512],prg3[2507:2504],prg3[2499:2496],
                  prg3[2491:2488],prg3[2483:2480],prg3[2475:2472],prg3[2467:2464],prg3[2459:2456],prg3[2451:2448],prg3[2443:2440],prg3[2435:2432],
                  prg3[2427:2424],prg3[2419:2416],prg3[2411:2408],prg3[2403:2400],prg3[2395:2392],prg3[2387:2384],prg3[2379:2376],prg3[2371:2368],
                  prg3[2363:2360],prg3[2355:2352],prg3[2347:2344],prg3[2339:2336],prg3[2331:2328],prg3[2323:2320],prg3[2315:2312],prg3[2307:2304],
                  prg3[2299:2296],prg3[2291:2288],prg3[2283:2280],prg3[2275:2272],prg3[2267:2264],prg3[2259:2256],prg3[2251:2248],prg3[2243:2240],
                  prg3[2235:2232],prg3[2227:2224],prg3[2219:2216],prg3[2211:2208],prg3[2203:2200],prg3[2195:2192],prg3[2187:2184],prg3[2179:2176],
                  prg3[2171:2168],prg3[2163:2160],prg3[2155:2152],prg3[2147:2144],prg3[2139:2136],prg3[2131:2128],prg3[2123:2120],prg3[2115:2112],
                  prg3[2107:2104],prg3[2099:2096],prg3[2091:2088],prg3[2083:2080],prg3[2075:2072],prg3[2067:2064],prg3[2059:2056],prg3[2051:2048],
                  prg3[2043:2040],prg3[2035:2032],prg3[2027:2024],prg3[2019:2016],prg3[2011:2008],prg3[2003:2000],prg3[1995:1992],prg3[1987:1984],
                  prg3[1979:1976],prg3[1971:1968],prg3[1963:1960],prg3[1955:1952],prg3[1947:1944],prg3[1939:1936],prg3[1931:1928],prg3[1923:1920],
                  prg3[1915:1912],prg3[1907:1904],prg3[1899:1896],prg3[1891:1888],prg3[1883:1880],prg3[1875:1872],prg3[1867:1864],prg3[1859:1856],
                  prg3[1851:1848],prg3[1843:1840],prg3[1835:1832],prg3[1827:1824],prg3[1819:1816],prg3[1811:1808],prg3[1803:1800],prg3[1795:1792],
                  prg3[1787:1784],prg3[1779:1776],prg3[1771:1768],prg3[1763:1760],prg3[1755:1752],prg3[1747:1744],prg3[1739:1736],prg3[1731:1728],
                  prg3[1723:1720],prg3[1715:1712],prg3[1707:1704],prg3[1699:1696],prg3[1691:1688],prg3[1683:1680],prg3[1675:1672],prg3[1667:1664],
                  prg3[1659:1656],prg3[1651:1648],prg3[1643:1640],prg3[1635:1632],prg3[1627:1624],prg3[1619:1616],prg3[1611:1608],prg3[1603:1600],
                  prg3[1595:1592],prg3[1587:1584],prg3[1579:1576],prg3[1571:1568],prg3[1563:1560],prg3[1555:1552],prg3[1547:1544],prg3[1539:1536],
                  prg3[1531:1528],prg3[1523:1520],prg3[1515:1512],prg3[1507:1504],prg3[1499:1496],prg3[1491:1488],prg3[1483:1480],prg3[1475:1472],
                  prg3[1467:1464],prg3[1459:1456],prg3[1451:1448],prg3[1443:1440],prg3[1435:1432],prg3[1427:1424],prg3[1419:1416],prg3[1411:1408],
                  prg3[1403:1400],prg3[1395:1392],prg3[1387:1384],prg3[1379:1376],prg3[1371:1368],prg3[1363:1360],prg3[1355:1352],prg3[1347:1344],
                  prg3[1339:1336],prg3[1331:1328],prg3[1323:1320],prg3[1315:1312],prg3[1307:1304],prg3[1299:1296],prg3[1291:1288],prg3[1283:1280],
                  prg3[1275:1272],prg3[1267:1264],prg3[1259:1256],prg3[1251:1248],prg3[1243:1240],prg3[1235:1232],prg3[1227:1224],prg3[1219:1216],
                  prg3[1211:1208],prg3[1203:1200],prg3[1195:1192],prg3[1187:1184],prg3[1179:1176],prg3[1171:1168],prg3[1163:1160],prg3[1155:1152],
                  prg3[1147:1144],prg3[1139:1136],prg3[1131:1128],prg3[1123:1120],prg3[1115:1112],prg3[1107:1104],prg3[1099:1096],prg3[1091:1088],
                  prg3[1083:1080],prg3[1075:1072],prg3[1067:1064],prg3[1059:1056],prg3[1051:1048],prg3[1043:1040],prg3[1035:1032],prg3[1027:1024],
                  prg3[1019:1016],prg3[1011:1008],prg3[1003:1000],prg3[ 995: 992],prg3[ 987: 984],prg3[ 979: 976],prg3[ 971: 968],prg3[ 963: 960],
                  prg3[ 955: 952],prg3[ 947: 944],prg3[ 939: 936],prg3[ 931: 928],prg3[ 923: 920],prg3[ 915: 912],prg3[ 907: 904],prg3[ 899: 896],
                  prg3[ 891: 888],prg3[ 883: 880],prg3[ 875: 872],prg3[ 867: 864],prg3[ 859: 856],prg3[ 851: 848],prg3[ 843: 840],prg3[ 835: 832],
                  prg3[ 827: 824],prg3[ 819: 816],prg3[ 811: 808],prg3[ 803: 800],prg3[ 795: 792],prg3[ 787: 784],prg3[ 779: 776],prg3[ 771: 768],
                  prg3[ 763: 760],prg3[ 755: 752],prg3[ 747: 744],prg3[ 739: 736],prg3[ 731: 728],prg3[ 723: 720],prg3[ 715: 712],prg3[ 707: 704],
                  prg3[ 699: 696],prg3[ 691: 688],prg3[ 683: 680],prg3[ 675: 672],prg3[ 667: 664],prg3[ 659: 656],prg3[ 651: 648],prg3[ 643: 640],
                  prg3[ 635: 632],prg3[ 627: 624],prg3[ 619: 616],prg3[ 611: 608],prg3[ 603: 600],prg3[ 595: 592],prg3[ 587: 584],prg3[ 579: 576],
                  prg3[ 571: 568],prg3[ 563: 560],prg3[ 555: 552],prg3[ 547: 544],prg3[ 539: 536],prg3[ 531: 528],prg3[ 523: 520],prg3[ 515: 512],
                  prg3[ 507: 504],prg3[ 499: 496],prg3[ 491: 488],prg3[ 483: 480],prg3[ 475: 472],prg3[ 467: 464],prg3[ 459: 456],prg3[ 451: 448],
                  prg3[ 443: 440],prg3[ 435: 432],prg3[ 427: 424],prg3[ 419: 416],prg3[ 411: 408],prg3[ 403: 400],prg3[ 395: 392],prg3[ 387: 384],
                  prg3[ 379: 376],prg3[ 371: 368],prg3[ 363: 360],prg3[ 355: 352],prg3[ 347: 344],prg3[ 339: 336],prg3[ 331: 328],prg3[ 323: 320],
                  prg3[ 315: 312],prg3[ 307: 304],prg3[ 299: 296],prg3[ 291: 288],prg3[ 283: 280],prg3[ 275: 272],prg3[ 267: 264],prg3[ 259: 256],
                  prg3[ 251: 248],prg3[ 243: 240],prg3[ 235: 232],prg3[ 227: 224],prg3[ 219: 216],prg3[ 211: 208],prg3[ 203: 200],prg3[ 195: 192],
                  prg3[ 187: 184],prg3[ 179: 176],prg3[ 171: 168],prg3[ 163: 160],prg3[ 155: 152],prg3[ 147: 144],prg3[ 139: 136],prg3[ 131: 128],
                  prg3[ 123: 120],prg3[ 115: 112],prg3[ 107: 104],prg3[  99:  96],prg3[  91:  88],prg3[  83:  80],prg3[  75:  72],prg3[  67:  64],
                  prg3[  59:  56],prg3[  51:  48],prg3[  43:  40],prg3[  35:  32],prg3[  27:  24],prg3[  19:  16],prg3[  11:   8],prg3[   3:   0],
                  prg2[4091:4088],prg2[4083:4080],prg2[4075:4072],prg2[4067:4064],prg2[4059:4056],prg2[4051:4048],prg2[4043:4040],prg2[4035:4032],
                  prg2[4027:4024],prg2[4019:4016],prg2[4011:4008],prg2[4003:4000],prg2[3995:3992],prg2[3987:3984],prg2[3979:3976],prg2[3971:3968],
                  prg2[3963:3960],prg2[3955:3952],prg2[3947:3944],prg2[3939:3936],prg2[3931:3928],prg2[3923:3920],prg2[3915:3912],prg2[3907:3904],
                  prg2[3899:3896],prg2[3891:3888],prg2[3883:3880],prg2[3875:3872],prg2[3867:3864],prg2[3859:3856],prg2[3851:3848],prg2[3843:3840],
                  prg2[3835:3832],prg2[3827:3824],prg2[3819:3816],prg2[3811:3808],prg2[3803:3800],prg2[3795:3792],prg2[3787:3784],prg2[3779:3776],
                  prg2[3771:3768],prg2[3763:3760],prg2[3755:3752],prg2[3747:3744],prg2[3739:3736],prg2[3731:3728],prg2[3723:3720],prg2[3715:3712],
                  prg2[3707:3704],prg2[3699:3696],prg2[3691:3688],prg2[3683:3680],prg2[3675:3672],prg2[3667:3664],prg2[3659:3656],prg2[3651:3648],
                  prg2[3643:3640],prg2[3635:3632],prg2[3627:3624],prg2[3619:3616],prg2[3611:3608],prg2[3603:3600],prg2[3595:3592],prg2[3587:3584],
                  prg2[3579:3576],prg2[3571:3568],prg2[3563:3560],prg2[3555:3552],prg2[3547:3544],prg2[3539:3536],prg2[3531:3528],prg2[3523:3520],
                  prg2[3515:3512],prg2[3507:3504],prg2[3499:3496],prg2[3491:3488],prg2[3483:3480],prg2[3475:3472],prg2[3467:3464],prg2[3459:3456],
                  prg2[3451:3448],prg2[3443:3440],prg2[3435:3432],prg2[3427:3424],prg2[3419:3416],prg2[3411:3408],prg2[3403:3400],prg2[3395:3392],
                  prg2[3387:3384],prg2[3379:3376],prg2[3371:3368],prg2[3363:3360],prg2[3355:3352],prg2[3347:3344],prg2[3339:3336],prg2[3331:3328],
                  prg2[3323:3320],prg2[3315:3312],prg2[3307:3304],prg2[3299:3296],prg2[3291:3288],prg2[3283:3280],prg2[3275:3272],prg2[3267:3264],
                  prg2[3259:3256],prg2[3251:3248],prg2[3243:3240],prg2[3235:3232],prg2[3227:3224],prg2[3219:3216],prg2[3211:3208],prg2[3203:3200],
                  prg2[3195:3192],prg2[3187:3184],prg2[3179:3176],prg2[3171:3168],prg2[3163:3160],prg2[3155:3152],prg2[3147:3144],prg2[3139:3136],
                  prg2[3131:3128],prg2[3123:3120],prg2[3115:3112],prg2[3107:3104],prg2[3099:3096],prg2[3091:3088],prg2[3083:3080],prg2[3075:3072],
                  prg2[3067:3064],prg2[3059:3056],prg2[3051:3048],prg2[3043:3040],prg2[3035:3032],prg2[3027:3024],prg2[3019:3016],prg2[3011:3008],
                  prg2[3003:3000],prg2[2995:2992],prg2[2987:2984],prg2[2979:2976],prg2[2971:2968],prg2[2963:2960],prg2[2955:2952],prg2[2947:2944],
                  prg2[2939:2936],prg2[2931:2928],prg2[2923:2920],prg2[2915:2912],prg2[2907:2904],prg2[2899:2896],prg2[2891:2888],prg2[2883:2880],
                  prg2[2875:2872],prg2[2867:2864],prg2[2859:2856],prg2[2851:2848],prg2[2843:2840],prg2[2835:2832],prg2[2827:2824],prg2[2819:2816],
                  prg2[2811:2808],prg2[2803:2800],prg2[2795:2792],prg2[2787:2784],prg2[2779:2776],prg2[2771:2768],prg2[2763:2760],prg2[2755:2752],
                  prg2[2747:2744],prg2[2739:2736],prg2[2731:2728],prg2[2723:2720],prg2[2715:2712],prg2[2707:2704],prg2[2699:2696],prg2[2691:2688],
                  prg2[2683:2680],prg2[2675:2672],prg2[2667:2664],prg2[2659:2656],prg2[2651:2648],prg2[2643:2640],prg2[2635:2632],prg2[2627:2624],
                  prg2[2619:2616],prg2[2611:2608],prg2[2603:2600],prg2[2595:2592],prg2[2587:2584],prg2[2579:2576],prg2[2571:2568],prg2[2563:2560],
                  prg2[2555:2552],prg2[2547:2544],prg2[2539:2536],prg2[2531:2528],prg2[2523:2520],prg2[2515:2512],prg2[2507:2504],prg2[2499:2496],
                  prg2[2491:2488],prg2[2483:2480],prg2[2475:2472],prg2[2467:2464],prg2[2459:2456],prg2[2451:2448],prg2[2443:2440],prg2[2435:2432],
                  prg2[2427:2424],prg2[2419:2416],prg2[2411:2408],prg2[2403:2400],prg2[2395:2392],prg2[2387:2384],prg2[2379:2376],prg2[2371:2368],
                  prg2[2363:2360],prg2[2355:2352],prg2[2347:2344],prg2[2339:2336],prg2[2331:2328],prg2[2323:2320],prg2[2315:2312],prg2[2307:2304],
                  prg2[2299:2296],prg2[2291:2288],prg2[2283:2280],prg2[2275:2272],prg2[2267:2264],prg2[2259:2256],prg2[2251:2248],prg2[2243:2240],
                  prg2[2235:2232],prg2[2227:2224],prg2[2219:2216],prg2[2211:2208],prg2[2203:2200],prg2[2195:2192],prg2[2187:2184],prg2[2179:2176],
                  prg2[2171:2168],prg2[2163:2160],prg2[2155:2152],prg2[2147:2144],prg2[2139:2136],prg2[2131:2128],prg2[2123:2120],prg2[2115:2112],
                  prg2[2107:2104],prg2[2099:2096],prg2[2091:2088],prg2[2083:2080],prg2[2075:2072],prg2[2067:2064],prg2[2059:2056],prg2[2051:2048],
                  prg2[2043:2040],prg2[2035:2032],prg2[2027:2024],prg2[2019:2016],prg2[2011:2008],prg2[2003:2000],prg2[1995:1992],prg2[1987:1984],
                  prg2[1979:1976],prg2[1971:1968],prg2[1963:1960],prg2[1955:1952],prg2[1947:1944],prg2[1939:1936],prg2[1931:1928],prg2[1923:1920],
                  prg2[1915:1912],prg2[1907:1904],prg2[1899:1896],prg2[1891:1888],prg2[1883:1880],prg2[1875:1872],prg2[1867:1864],prg2[1859:1856],
                  prg2[1851:1848],prg2[1843:1840],prg2[1835:1832],prg2[1827:1824],prg2[1819:1816],prg2[1811:1808],prg2[1803:1800],prg2[1795:1792],
                  prg2[1787:1784],prg2[1779:1776],prg2[1771:1768],prg2[1763:1760],prg2[1755:1752],prg2[1747:1744],prg2[1739:1736],prg2[1731:1728],
                  prg2[1723:1720],prg2[1715:1712],prg2[1707:1704],prg2[1699:1696],prg2[1691:1688],prg2[1683:1680],prg2[1675:1672],prg2[1667:1664],
                  prg2[1659:1656],prg2[1651:1648],prg2[1643:1640],prg2[1635:1632],prg2[1627:1624],prg2[1619:1616],prg2[1611:1608],prg2[1603:1600],
                  prg2[1595:1592],prg2[1587:1584],prg2[1579:1576],prg2[1571:1568],prg2[1563:1560],prg2[1555:1552],prg2[1547:1544],prg2[1539:1536],
                  prg2[1531:1528],prg2[1523:1520],prg2[1515:1512],prg2[1507:1504],prg2[1499:1496],prg2[1491:1488],prg2[1483:1480],prg2[1475:1472],
                  prg2[1467:1464],prg2[1459:1456],prg2[1451:1448],prg2[1443:1440],prg2[1435:1432],prg2[1427:1424],prg2[1419:1416],prg2[1411:1408],
                  prg2[1403:1400],prg2[1395:1392],prg2[1387:1384],prg2[1379:1376],prg2[1371:1368],prg2[1363:1360],prg2[1355:1352],prg2[1347:1344],
                  prg2[1339:1336],prg2[1331:1328],prg2[1323:1320],prg2[1315:1312],prg2[1307:1304],prg2[1299:1296],prg2[1291:1288],prg2[1283:1280],
                  prg2[1275:1272],prg2[1267:1264],prg2[1259:1256],prg2[1251:1248],prg2[1243:1240],prg2[1235:1232],prg2[1227:1224],prg2[1219:1216],
                  prg2[1211:1208],prg2[1203:1200],prg2[1195:1192],prg2[1187:1184],prg2[1179:1176],prg2[1171:1168],prg2[1163:1160],prg2[1155:1152],
                  prg2[1147:1144],prg2[1139:1136],prg2[1131:1128],prg2[1123:1120],prg2[1115:1112],prg2[1107:1104],prg2[1099:1096],prg2[1091:1088],
                  prg2[1083:1080],prg2[1075:1072],prg2[1067:1064],prg2[1059:1056],prg2[1051:1048],prg2[1043:1040],prg2[1035:1032],prg2[1027:1024],
                  prg2[1019:1016],prg2[1011:1008],prg2[1003:1000],prg2[ 995: 992],prg2[ 987: 984],prg2[ 979: 976],prg2[ 971: 968],prg2[ 963: 960],
                  prg2[ 955: 952],prg2[ 947: 944],prg2[ 939: 936],prg2[ 931: 928],prg2[ 923: 920],prg2[ 915: 912],prg2[ 907: 904],prg2[ 899: 896],
                  prg2[ 891: 888],prg2[ 883: 880],prg2[ 875: 872],prg2[ 867: 864],prg2[ 859: 856],prg2[ 851: 848],prg2[ 843: 840],prg2[ 835: 832],
                  prg2[ 827: 824],prg2[ 819: 816],prg2[ 811: 808],prg2[ 803: 800],prg2[ 795: 792],prg2[ 787: 784],prg2[ 779: 776],prg2[ 771: 768],
                  prg2[ 763: 760],prg2[ 755: 752],prg2[ 747: 744],prg2[ 739: 736],prg2[ 731: 728],prg2[ 723: 720],prg2[ 715: 712],prg2[ 707: 704],
                  prg2[ 699: 696],prg2[ 691: 688],prg2[ 683: 680],prg2[ 675: 672],prg2[ 667: 664],prg2[ 659: 656],prg2[ 651: 648],prg2[ 643: 640],
                  prg2[ 635: 632],prg2[ 627: 624],prg2[ 619: 616],prg2[ 611: 608],prg2[ 603: 600],prg2[ 595: 592],prg2[ 587: 584],prg2[ 579: 576],
                  prg2[ 571: 568],prg2[ 563: 560],prg2[ 555: 552],prg2[ 547: 544],prg2[ 539: 536],prg2[ 531: 528],prg2[ 523: 520],prg2[ 515: 512],
                  prg2[ 507: 504],prg2[ 499: 496],prg2[ 491: 488],prg2[ 483: 480],prg2[ 475: 472],prg2[ 467: 464],prg2[ 459: 456],prg2[ 451: 448],
                  prg2[ 443: 440],prg2[ 435: 432],prg2[ 427: 424],prg2[ 419: 416],prg2[ 411: 408],prg2[ 403: 400],prg2[ 395: 392],prg2[ 387: 384],
                  prg2[ 379: 376],prg2[ 371: 368],prg2[ 363: 360],prg2[ 355: 352],prg2[ 347: 344],prg2[ 339: 336],prg2[ 331: 328],prg2[ 323: 320],
                  prg2[ 315: 312],prg2[ 307: 304],prg2[ 299: 296],prg2[ 291: 288],prg2[ 283: 280],prg2[ 275: 272],prg2[ 267: 264],prg2[ 259: 256],
                  prg2[ 251: 248],prg2[ 243: 240],prg2[ 235: 232],prg2[ 227: 224],prg2[ 219: 216],prg2[ 211: 208],prg2[ 203: 200],prg2[ 195: 192],
                  prg2[ 187: 184],prg2[ 179: 176],prg2[ 171: 168],prg2[ 163: 160],prg2[ 155: 152],prg2[ 147: 144],prg2[ 139: 136],prg2[ 131: 128],
                  prg2[ 123: 120],prg2[ 115: 112],prg2[ 107: 104],prg2[  99:  96],prg2[  91:  88],prg2[  83:  80],prg2[  75:  72],prg2[  67:  64],
                  prg2[  59:  56],prg2[  51:  48],prg2[  43:  40],prg2[  35:  32],prg2[  27:  24],prg2[  19:  16],prg2[  11:   8],prg2[   3:   0]};
         localparam [4095:0]
           pb0 = {prg1[4091:4088],prg1[4083:4080],prg1[4075:4072],prg1[4067:4064],prg1[4059:4056],prg1[4051:4048],prg1[4043:4040],prg1[4035:4032],
                  prg1[4027:4024],prg1[4019:4016],prg1[4011:4008],prg1[4003:4000],prg1[3995:3992],prg1[3987:3984],prg1[3979:3976],prg1[3971:3968],
                  prg1[3963:3960],prg1[3955:3952],prg1[3947:3944],prg1[3939:3936],prg1[3931:3928],prg1[3923:3920],prg1[3915:3912],prg1[3907:3904],
                  prg1[3899:3896],prg1[3891:3888],prg1[3883:3880],prg1[3875:3872],prg1[3867:3864],prg1[3859:3856],prg1[3851:3848],prg1[3843:3840],
                  prg1[3835:3832],prg1[3827:3824],prg1[3819:3816],prg1[3811:3808],prg1[3803:3800],prg1[3795:3792],prg1[3787:3784],prg1[3779:3776],
                  prg1[3771:3768],prg1[3763:3760],prg1[3755:3752],prg1[3747:3744],prg1[3739:3736],prg1[3731:3728],prg1[3723:3720],prg1[3715:3712],
                  prg1[3707:3704],prg1[3699:3696],prg1[3691:3688],prg1[3683:3680],prg1[3675:3672],prg1[3667:3664],prg1[3659:3656],prg1[3651:3648],
                  prg1[3643:3640],prg1[3635:3632],prg1[3627:3624],prg1[3619:3616],prg1[3611:3608],prg1[3603:3600],prg1[3595:3592],prg1[3587:3584],
                  prg1[3579:3576],prg1[3571:3568],prg1[3563:3560],prg1[3555:3552],prg1[3547:3544],prg1[3539:3536],prg1[3531:3528],prg1[3523:3520],
                  prg1[3515:3512],prg1[3507:3504],prg1[3499:3496],prg1[3491:3488],prg1[3483:3480],prg1[3475:3472],prg1[3467:3464],prg1[3459:3456],
                  prg1[3451:3448],prg1[3443:3440],prg1[3435:3432],prg1[3427:3424],prg1[3419:3416],prg1[3411:3408],prg1[3403:3400],prg1[3395:3392],
                  prg1[3387:3384],prg1[3379:3376],prg1[3371:3368],prg1[3363:3360],prg1[3355:3352],prg1[3347:3344],prg1[3339:3336],prg1[3331:3328],
                  prg1[3323:3320],prg1[3315:3312],prg1[3307:3304],prg1[3299:3296],prg1[3291:3288],prg1[3283:3280],prg1[3275:3272],prg1[3267:3264],
                  prg1[3259:3256],prg1[3251:3248],prg1[3243:3240],prg1[3235:3232],prg1[3227:3224],prg1[3219:3216],prg1[3211:3208],prg1[3203:3200],
                  prg1[3195:3192],prg1[3187:3184],prg1[3179:3176],prg1[3171:3168],prg1[3163:3160],prg1[3155:3152],prg1[3147:3144],prg1[3139:3136],
                  prg1[3131:3128],prg1[3123:3120],prg1[3115:3112],prg1[3107:3104],prg1[3099:3096],prg1[3091:3088],prg1[3083:3080],prg1[3075:3072],
                  prg1[3067:3064],prg1[3059:3056],prg1[3051:3048],prg1[3043:3040],prg1[3035:3032],prg1[3027:3024],prg1[3019:3016],prg1[3011:3008],
                  prg1[3003:3000],prg1[2995:2992],prg1[2987:2984],prg1[2979:2976],prg1[2971:2968],prg1[2963:2960],prg1[2955:2952],prg1[2947:2944],
                  prg1[2939:2936],prg1[2931:2928],prg1[2923:2920],prg1[2915:2912],prg1[2907:2904],prg1[2899:2896],prg1[2891:2888],prg1[2883:2880],
                  prg1[2875:2872],prg1[2867:2864],prg1[2859:2856],prg1[2851:2848],prg1[2843:2840],prg1[2835:2832],prg1[2827:2824],prg1[2819:2816],
                  prg1[2811:2808],prg1[2803:2800],prg1[2795:2792],prg1[2787:2784],prg1[2779:2776],prg1[2771:2768],prg1[2763:2760],prg1[2755:2752],
                  prg1[2747:2744],prg1[2739:2736],prg1[2731:2728],prg1[2723:2720],prg1[2715:2712],prg1[2707:2704],prg1[2699:2696],prg1[2691:2688],
                  prg1[2683:2680],prg1[2675:2672],prg1[2667:2664],prg1[2659:2656],prg1[2651:2648],prg1[2643:2640],prg1[2635:2632],prg1[2627:2624],
                  prg1[2619:2616],prg1[2611:2608],prg1[2603:2600],prg1[2595:2592],prg1[2587:2584],prg1[2579:2576],prg1[2571:2568],prg1[2563:2560],
                  prg1[2555:2552],prg1[2547:2544],prg1[2539:2536],prg1[2531:2528],prg1[2523:2520],prg1[2515:2512],prg1[2507:2504],prg1[2499:2496],
                  prg1[2491:2488],prg1[2483:2480],prg1[2475:2472],prg1[2467:2464],prg1[2459:2456],prg1[2451:2448],prg1[2443:2440],prg1[2435:2432],
                  prg1[2427:2424],prg1[2419:2416],prg1[2411:2408],prg1[2403:2400],prg1[2395:2392],prg1[2387:2384],prg1[2379:2376],prg1[2371:2368],
                  prg1[2363:2360],prg1[2355:2352],prg1[2347:2344],prg1[2339:2336],prg1[2331:2328],prg1[2323:2320],prg1[2315:2312],prg1[2307:2304],
                  prg1[2299:2296],prg1[2291:2288],prg1[2283:2280],prg1[2275:2272],prg1[2267:2264],prg1[2259:2256],prg1[2251:2248],prg1[2243:2240],
                  prg1[2235:2232],prg1[2227:2224],prg1[2219:2216],prg1[2211:2208],prg1[2203:2200],prg1[2195:2192],prg1[2187:2184],prg1[2179:2176],
                  prg1[2171:2168],prg1[2163:2160],prg1[2155:2152],prg1[2147:2144],prg1[2139:2136],prg1[2131:2128],prg1[2123:2120],prg1[2115:2112],
                  prg1[2107:2104],prg1[2099:2096],prg1[2091:2088],prg1[2083:2080],prg1[2075:2072],prg1[2067:2064],prg1[2059:2056],prg1[2051:2048],
                  prg1[2043:2040],prg1[2035:2032],prg1[2027:2024],prg1[2019:2016],prg1[2011:2008],prg1[2003:2000],prg1[1995:1992],prg1[1987:1984],
                  prg1[1979:1976],prg1[1971:1968],prg1[1963:1960],prg1[1955:1952],prg1[1947:1944],prg1[1939:1936],prg1[1931:1928],prg1[1923:1920],
                  prg1[1915:1912],prg1[1907:1904],prg1[1899:1896],prg1[1891:1888],prg1[1883:1880],prg1[1875:1872],prg1[1867:1864],prg1[1859:1856],
                  prg1[1851:1848],prg1[1843:1840],prg1[1835:1832],prg1[1827:1824],prg1[1819:1816],prg1[1811:1808],prg1[1803:1800],prg1[1795:1792],
                  prg1[1787:1784],prg1[1779:1776],prg1[1771:1768],prg1[1763:1760],prg1[1755:1752],prg1[1747:1744],prg1[1739:1736],prg1[1731:1728],
                  prg1[1723:1720],prg1[1715:1712],prg1[1707:1704],prg1[1699:1696],prg1[1691:1688],prg1[1683:1680],prg1[1675:1672],prg1[1667:1664],
                  prg1[1659:1656],prg1[1651:1648],prg1[1643:1640],prg1[1635:1632],prg1[1627:1624],prg1[1619:1616],prg1[1611:1608],prg1[1603:1600],
                  prg1[1595:1592],prg1[1587:1584],prg1[1579:1576],prg1[1571:1568],prg1[1563:1560],prg1[1555:1552],prg1[1547:1544],prg1[1539:1536],
                  prg1[1531:1528],prg1[1523:1520],prg1[1515:1512],prg1[1507:1504],prg1[1499:1496],prg1[1491:1488],prg1[1483:1480],prg1[1475:1472],
                  prg1[1467:1464],prg1[1459:1456],prg1[1451:1448],prg1[1443:1440],prg1[1435:1432],prg1[1427:1424],prg1[1419:1416],prg1[1411:1408],
                  prg1[1403:1400],prg1[1395:1392],prg1[1387:1384],prg1[1379:1376],prg1[1371:1368],prg1[1363:1360],prg1[1355:1352],prg1[1347:1344],
                  prg1[1339:1336],prg1[1331:1328],prg1[1323:1320],prg1[1315:1312],prg1[1307:1304],prg1[1299:1296],prg1[1291:1288],prg1[1283:1280],
                  prg1[1275:1272],prg1[1267:1264],prg1[1259:1256],prg1[1251:1248],prg1[1243:1240],prg1[1235:1232],prg1[1227:1224],prg1[1219:1216],
                  prg1[1211:1208],prg1[1203:1200],prg1[1195:1192],prg1[1187:1184],prg1[1179:1176],prg1[1171:1168],prg1[1163:1160],prg1[1155:1152],
                  prg1[1147:1144],prg1[1139:1136],prg1[1131:1128],prg1[1123:1120],prg1[1115:1112],prg1[1107:1104],prg1[1099:1096],prg1[1091:1088],
                  prg1[1083:1080],prg1[1075:1072],prg1[1067:1064],prg1[1059:1056],prg1[1051:1048],prg1[1043:1040],prg1[1035:1032],prg1[1027:1024],
                  prg1[1019:1016],prg1[1011:1008],prg1[1003:1000],prg1[ 995: 992],prg1[ 987: 984],prg1[ 979: 976],prg1[ 971: 968],prg1[ 963: 960],
                  prg1[ 955: 952],prg1[ 947: 944],prg1[ 939: 936],prg1[ 931: 928],prg1[ 923: 920],prg1[ 915: 912],prg1[ 907: 904],prg1[ 899: 896],
                  prg1[ 891: 888],prg1[ 883: 880],prg1[ 875: 872],prg1[ 867: 864],prg1[ 859: 856],prg1[ 851: 848],prg1[ 843: 840],prg1[ 835: 832],
                  prg1[ 827: 824],prg1[ 819: 816],prg1[ 811: 808],prg1[ 803: 800],prg1[ 795: 792],prg1[ 787: 784],prg1[ 779: 776],prg1[ 771: 768],
                  prg1[ 763: 760],prg1[ 755: 752],prg1[ 747: 744],prg1[ 739: 736],prg1[ 731: 728],prg1[ 723: 720],prg1[ 715: 712],prg1[ 707: 704],
                  prg1[ 699: 696],prg1[ 691: 688],prg1[ 683: 680],prg1[ 675: 672],prg1[ 667: 664],prg1[ 659: 656],prg1[ 651: 648],prg1[ 643: 640],
                  prg1[ 635: 632],prg1[ 627: 624],prg1[ 619: 616],prg1[ 611: 608],prg1[ 603: 600],prg1[ 595: 592],prg1[ 587: 584],prg1[ 579: 576],
                  prg1[ 571: 568],prg1[ 563: 560],prg1[ 555: 552],prg1[ 547: 544],prg1[ 539: 536],prg1[ 531: 528],prg1[ 523: 520],prg1[ 515: 512],
                  prg1[ 507: 504],prg1[ 499: 496],prg1[ 491: 488],prg1[ 483: 480],prg1[ 475: 472],prg1[ 467: 464],prg1[ 459: 456],prg1[ 451: 448],
                  prg1[ 443: 440],prg1[ 435: 432],prg1[ 427: 424],prg1[ 419: 416],prg1[ 411: 408],prg1[ 403: 400],prg1[ 395: 392],prg1[ 387: 384],
                  prg1[ 379: 376],prg1[ 371: 368],prg1[ 363: 360],prg1[ 355: 352],prg1[ 347: 344],prg1[ 339: 336],prg1[ 331: 328],prg1[ 323: 320],
                  prg1[ 315: 312],prg1[ 307: 304],prg1[ 299: 296],prg1[ 291: 288],prg1[ 283: 280],prg1[ 275: 272],prg1[ 267: 264],prg1[ 259: 256],
                  prg1[ 251: 248],prg1[ 243: 240],prg1[ 235: 232],prg1[ 227: 224],prg1[ 219: 216],prg1[ 211: 208],prg1[ 203: 200],prg1[ 195: 192],
                  prg1[ 187: 184],prg1[ 179: 176],prg1[ 171: 168],prg1[ 163: 160],prg1[ 155: 152],prg1[ 147: 144],prg1[ 139: 136],prg1[ 131: 128],
                  prg1[ 123: 120],prg1[ 115: 112],prg1[ 107: 104],prg1[  99:  96],prg1[  91:  88],prg1[  83:  80],prg1[  75:  72],prg1[  67:  64],
                  prg1[  59:  56],prg1[  51:  48],prg1[  43:  40],prg1[  35:  32],prg1[  27:  24],prg1[  19:  16],prg1[  11:   8],prg1[   3:   0],
                  prg0[4091:4088],prg0[4083:4080],prg0[4075:4072],prg0[4067:4064],prg0[4059:4056],prg0[4051:4048],prg0[4043:4040],prg0[4035:4032],
                  prg0[4027:4024],prg0[4019:4016],prg0[4011:4008],prg0[4003:4000],prg0[3995:3992],prg0[3987:3984],prg0[3979:3976],prg0[3971:3968],
                  prg0[3963:3960],prg0[3955:3952],prg0[3947:3944],prg0[3939:3936],prg0[3931:3928],prg0[3923:3920],prg0[3915:3912],prg0[3907:3904],
                  prg0[3899:3896],prg0[3891:3888],prg0[3883:3880],prg0[3875:3872],prg0[3867:3864],prg0[3859:3856],prg0[3851:3848],prg0[3843:3840],
                  prg0[3835:3832],prg0[3827:3824],prg0[3819:3816],prg0[3811:3808],prg0[3803:3800],prg0[3795:3792],prg0[3787:3784],prg0[3779:3776],
                  prg0[3771:3768],prg0[3763:3760],prg0[3755:3752],prg0[3747:3744],prg0[3739:3736],prg0[3731:3728],prg0[3723:3720],prg0[3715:3712],
                  prg0[3707:3704],prg0[3699:3696],prg0[3691:3688],prg0[3683:3680],prg0[3675:3672],prg0[3667:3664],prg0[3659:3656],prg0[3651:3648],
                  prg0[3643:3640],prg0[3635:3632],prg0[3627:3624],prg0[3619:3616],prg0[3611:3608],prg0[3603:3600],prg0[3595:3592],prg0[3587:3584],
                  prg0[3579:3576],prg0[3571:3568],prg0[3563:3560],prg0[3555:3552],prg0[3547:3544],prg0[3539:3536],prg0[3531:3528],prg0[3523:3520],
                  prg0[3515:3512],prg0[3507:3504],prg0[3499:3496],prg0[3491:3488],prg0[3483:3480],prg0[3475:3472],prg0[3467:3464],prg0[3459:3456],
                  prg0[3451:3448],prg0[3443:3440],prg0[3435:3432],prg0[3427:3424],prg0[3419:3416],prg0[3411:3408],prg0[3403:3400],prg0[3395:3392],
                  prg0[3387:3384],prg0[3379:3376],prg0[3371:3368],prg0[3363:3360],prg0[3355:3352],prg0[3347:3344],prg0[3339:3336],prg0[3331:3328],
                  prg0[3323:3320],prg0[3315:3312],prg0[3307:3304],prg0[3299:3296],prg0[3291:3288],prg0[3283:3280],prg0[3275:3272],prg0[3267:3264],
                  prg0[3259:3256],prg0[3251:3248],prg0[3243:3240],prg0[3235:3232],prg0[3227:3224],prg0[3219:3216],prg0[3211:3208],prg0[3203:3200],
                  prg0[3195:3192],prg0[3187:3184],prg0[3179:3176],prg0[3171:3168],prg0[3163:3160],prg0[3155:3152],prg0[3147:3144],prg0[3139:3136],
                  prg0[3131:3128],prg0[3123:3120],prg0[3115:3112],prg0[3107:3104],prg0[3099:3096],prg0[3091:3088],prg0[3083:3080],prg0[3075:3072],
                  prg0[3067:3064],prg0[3059:3056],prg0[3051:3048],prg0[3043:3040],prg0[3035:3032],prg0[3027:3024],prg0[3019:3016],prg0[3011:3008],
                  prg0[3003:3000],prg0[2995:2992],prg0[2987:2984],prg0[2979:2976],prg0[2971:2968],prg0[2963:2960],prg0[2955:2952],prg0[2947:2944],
                  prg0[2939:2936],prg0[2931:2928],prg0[2923:2920],prg0[2915:2912],prg0[2907:2904],prg0[2899:2896],prg0[2891:2888],prg0[2883:2880],
                  prg0[2875:2872],prg0[2867:2864],prg0[2859:2856],prg0[2851:2848],prg0[2843:2840],prg0[2835:2832],prg0[2827:2824],prg0[2819:2816],
                  prg0[2811:2808],prg0[2803:2800],prg0[2795:2792],prg0[2787:2784],prg0[2779:2776],prg0[2771:2768],prg0[2763:2760],prg0[2755:2752],
                  prg0[2747:2744],prg0[2739:2736],prg0[2731:2728],prg0[2723:2720],prg0[2715:2712],prg0[2707:2704],prg0[2699:2696],prg0[2691:2688],
                  prg0[2683:2680],prg0[2675:2672],prg0[2667:2664],prg0[2659:2656],prg0[2651:2648],prg0[2643:2640],prg0[2635:2632],prg0[2627:2624],
                  prg0[2619:2616],prg0[2611:2608],prg0[2603:2600],prg0[2595:2592],prg0[2587:2584],prg0[2579:2576],prg0[2571:2568],prg0[2563:2560],
                  prg0[2555:2552],prg0[2547:2544],prg0[2539:2536],prg0[2531:2528],prg0[2523:2520],prg0[2515:2512],prg0[2507:2504],prg0[2499:2496],
                  prg0[2491:2488],prg0[2483:2480],prg0[2475:2472],prg0[2467:2464],prg0[2459:2456],prg0[2451:2448],prg0[2443:2440],prg0[2435:2432],
                  prg0[2427:2424],prg0[2419:2416],prg0[2411:2408],prg0[2403:2400],prg0[2395:2392],prg0[2387:2384],prg0[2379:2376],prg0[2371:2368],
                  prg0[2363:2360],prg0[2355:2352],prg0[2347:2344],prg0[2339:2336],prg0[2331:2328],prg0[2323:2320],prg0[2315:2312],prg0[2307:2304],
                  prg0[2299:2296],prg0[2291:2288],prg0[2283:2280],prg0[2275:2272],prg0[2267:2264],prg0[2259:2256],prg0[2251:2248],prg0[2243:2240],
                  prg0[2235:2232],prg0[2227:2224],prg0[2219:2216],prg0[2211:2208],prg0[2203:2200],prg0[2195:2192],prg0[2187:2184],prg0[2179:2176],
                  prg0[2171:2168],prg0[2163:2160],prg0[2155:2152],prg0[2147:2144],prg0[2139:2136],prg0[2131:2128],prg0[2123:2120],prg0[2115:2112],
                  prg0[2107:2104],prg0[2099:2096],prg0[2091:2088],prg0[2083:2080],prg0[2075:2072],prg0[2067:2064],prg0[2059:2056],prg0[2051:2048],
                  prg0[2043:2040],prg0[2035:2032],prg0[2027:2024],prg0[2019:2016],prg0[2011:2008],prg0[2003:2000],prg0[1995:1992],prg0[1987:1984],
                  prg0[1979:1976],prg0[1971:1968],prg0[1963:1960],prg0[1955:1952],prg0[1947:1944],prg0[1939:1936],prg0[1931:1928],prg0[1923:1920],
                  prg0[1915:1912],prg0[1907:1904],prg0[1899:1896],prg0[1891:1888],prg0[1883:1880],prg0[1875:1872],prg0[1867:1864],prg0[1859:1856],
                  prg0[1851:1848],prg0[1843:1840],prg0[1835:1832],prg0[1827:1824],prg0[1819:1816],prg0[1811:1808],prg0[1803:1800],prg0[1795:1792],
                  prg0[1787:1784],prg0[1779:1776],prg0[1771:1768],prg0[1763:1760],prg0[1755:1752],prg0[1747:1744],prg0[1739:1736],prg0[1731:1728],
                  prg0[1723:1720],prg0[1715:1712],prg0[1707:1704],prg0[1699:1696],prg0[1691:1688],prg0[1683:1680],prg0[1675:1672],prg0[1667:1664],
                  prg0[1659:1656],prg0[1651:1648],prg0[1643:1640],prg0[1635:1632],prg0[1627:1624],prg0[1619:1616],prg0[1611:1608],prg0[1603:1600],
                  prg0[1595:1592],prg0[1587:1584],prg0[1579:1576],prg0[1571:1568],prg0[1563:1560],prg0[1555:1552],prg0[1547:1544],prg0[1539:1536],
                  prg0[1531:1528],prg0[1523:1520],prg0[1515:1512],prg0[1507:1504],prg0[1499:1496],prg0[1491:1488],prg0[1483:1480],prg0[1475:1472],
                  prg0[1467:1464],prg0[1459:1456],prg0[1451:1448],prg0[1443:1440],prg0[1435:1432],prg0[1427:1424],prg0[1419:1416],prg0[1411:1408],
                  prg0[1403:1400],prg0[1395:1392],prg0[1387:1384],prg0[1379:1376],prg0[1371:1368],prg0[1363:1360],prg0[1355:1352],prg0[1347:1344],
                  prg0[1339:1336],prg0[1331:1328],prg0[1323:1320],prg0[1315:1312],prg0[1307:1304],prg0[1299:1296],prg0[1291:1288],prg0[1283:1280],
                  prg0[1275:1272],prg0[1267:1264],prg0[1259:1256],prg0[1251:1248],prg0[1243:1240],prg0[1235:1232],prg0[1227:1224],prg0[1219:1216],
                  prg0[1211:1208],prg0[1203:1200],prg0[1195:1192],prg0[1187:1184],prg0[1179:1176],prg0[1171:1168],prg0[1163:1160],prg0[1155:1152],
                  prg0[1147:1144],prg0[1139:1136],prg0[1131:1128],prg0[1123:1120],prg0[1115:1112],prg0[1107:1104],prg0[1099:1096],prg0[1091:1088],
                  prg0[1083:1080],prg0[1075:1072],prg0[1067:1064],prg0[1059:1056],prg0[1051:1048],prg0[1043:1040],prg0[1035:1032],prg0[1027:1024],
                  prg0[1019:1016],prg0[1011:1008],prg0[1003:1000],prg0[ 995: 992],prg0[ 987: 984],prg0[ 979: 976],prg0[ 971: 968],prg0[ 963: 960],
                  prg0[ 955: 952],prg0[ 947: 944],prg0[ 939: 936],prg0[ 931: 928],prg0[ 923: 920],prg0[ 915: 912],prg0[ 907: 904],prg0[ 899: 896],
                  prg0[ 891: 888],prg0[ 883: 880],prg0[ 875: 872],prg0[ 867: 864],prg0[ 859: 856],prg0[ 851: 848],prg0[ 843: 840],prg0[ 835: 832],
                  prg0[ 827: 824],prg0[ 819: 816],prg0[ 811: 808],prg0[ 803: 800],prg0[ 795: 792],prg0[ 787: 784],prg0[ 779: 776],prg0[ 771: 768],
                  prg0[ 763: 760],prg0[ 755: 752],prg0[ 747: 744],prg0[ 739: 736],prg0[ 731: 728],prg0[ 723: 720],prg0[ 715: 712],prg0[ 707: 704],
                  prg0[ 699: 696],prg0[ 691: 688],prg0[ 683: 680],prg0[ 675: 672],prg0[ 667: 664],prg0[ 659: 656],prg0[ 651: 648],prg0[ 643: 640],
                  prg0[ 635: 632],prg0[ 627: 624],prg0[ 619: 616],prg0[ 611: 608],prg0[ 603: 600],prg0[ 595: 592],prg0[ 587: 584],prg0[ 579: 576],
                  prg0[ 571: 568],prg0[ 563: 560],prg0[ 555: 552],prg0[ 547: 544],prg0[ 539: 536],prg0[ 531: 528],prg0[ 523: 520],prg0[ 515: 512],
                  prg0[ 507: 504],prg0[ 499: 496],prg0[ 491: 488],prg0[ 483: 480],prg0[ 475: 472],prg0[ 467: 464],prg0[ 459: 456],prg0[ 451: 448],
                  prg0[ 443: 440],prg0[ 435: 432],prg0[ 427: 424],prg0[ 419: 416],prg0[ 411: 408],prg0[ 403: 400],prg0[ 395: 392],prg0[ 387: 384],
                  prg0[ 379: 376],prg0[ 371: 368],prg0[ 363: 360],prg0[ 355: 352],prg0[ 347: 344],prg0[ 339: 336],prg0[ 331: 328],prg0[ 323: 320],
                  prg0[ 315: 312],prg0[ 307: 304],prg0[ 299: 296],prg0[ 291: 288],prg0[ 283: 280],prg0[ 275: 272],prg0[ 267: 264],prg0[ 259: 256],
                  prg0[ 251: 248],prg0[ 243: 240],prg0[ 235: 232],prg0[ 227: 224],prg0[ 219: 216],prg0[ 211: 208],prg0[ 203: 200],prg0[ 195: 192],
                  prg0[ 187: 184],prg0[ 179: 176],prg0[ 171: 168],prg0[ 163: 160],prg0[ 155: 152],prg0[ 147: 144],prg0[ 139: 136],prg0[ 131: 128],
                  prg0[ 123: 120],prg0[ 115: 112],prg0[ 107: 104],prg0[  99:  96],prg0[  91:  88],prg0[  83:  80],prg0[  75:  72],prg0[  67:  64],
                  prg0[  59:  56],prg0[  51:  48],prg0[  43:  40],prg0[  35:  32],prg0[  27:  24],prg0[  19:  16],prg0[  11:   8],prg0[   3:   0]};
         localparam [4095:0]
           ph1 = {prg3[4095:4092],prg3[4087:4084],prg3[4079:4076],prg3[4071:4068],prg3[4063:4060],prg3[4055:4052],prg3[4047:4044],prg3[4039:4036],
                  prg3[4031:4028],prg3[4023:4020],prg3[4015:4012],prg3[4007:4004],prg3[3999:3996],prg3[3991:3988],prg3[3983:3980],prg3[3975:3972],
                  prg3[3967:3964],prg3[3959:3956],prg3[3951:3948],prg3[3943:3940],prg3[3935:3932],prg3[3927:3924],prg3[3919:3916],prg3[3911:3908],
                  prg3[3903:3900],prg3[3895:3892],prg3[3887:3884],prg3[3879:3876],prg3[3871:3868],prg3[3863:3860],prg3[3855:3852],prg3[3847:3844],
                  prg3[3839:3836],prg3[3831:3828],prg3[3823:3820],prg3[3815:3812],prg3[3807:3804],prg3[3799:3796],prg3[3791:3788],prg3[3783:3780],
                  prg3[3775:3772],prg3[3767:3764],prg3[3759:3756],prg3[3751:3748],prg3[3743:3740],prg3[3735:3732],prg3[3727:3724],prg3[3719:3716],
                  prg3[3711:3708],prg3[3703:3700],prg3[3695:3692],prg3[3687:3684],prg3[3679:3676],prg3[3671:3668],prg3[3663:3660],prg3[3655:3652],
                  prg3[3647:3644],prg3[3639:3636],prg3[3631:3628],prg3[3623:3620],prg3[3615:3612],prg3[3607:3604],prg3[3599:3596],prg3[3591:3588],
                  prg3[3583:3580],prg3[3575:3572],prg3[3567:3564],prg3[3559:3556],prg3[3551:3548],prg3[3543:3540],prg3[3535:3532],prg3[3527:3524],
                  prg3[3519:3516],prg3[3511:3508],prg3[3503:3500],prg3[3495:3492],prg3[3487:3484],prg3[3479:3476],prg3[3471:3468],prg3[3463:3460],
                  prg3[3455:3452],prg3[3447:3444],prg3[3439:3436],prg3[3431:3428],prg3[3423:3420],prg3[3415:3412],prg3[3407:3404],prg3[3399:3396],
                  prg3[3391:3388],prg3[3383:3380],prg3[3375:3372],prg3[3367:3364],prg3[3359:3356],prg3[3351:3348],prg3[3343:3340],prg3[3335:3332],
                  prg3[3327:3324],prg3[3319:3316],prg3[3311:3308],prg3[3303:3300],prg3[3295:3292],prg3[3287:3284],prg3[3279:3276],prg3[3271:3268],
                  prg3[3263:3260],prg3[3255:3252],prg3[3247:3244],prg3[3239:3236],prg3[3231:3228],prg3[3223:3220],prg3[3215:3212],prg3[3207:3204],
                  prg3[3199:3196],prg3[3191:3188],prg3[3183:3180],prg3[3175:3172],prg3[3167:3164],prg3[3159:3156],prg3[3151:3148],prg3[3143:3140],
                  prg3[3135:3132],prg3[3127:3124],prg3[3119:3116],prg3[3111:3108],prg3[3103:3100],prg3[3095:3092],prg3[3087:3084],prg3[3079:3076],
                  prg3[3071:3068],prg3[3063:3060],prg3[3055:3052],prg3[3047:3044],prg3[3039:3036],prg3[3031:3028],prg3[3023:3020],prg3[3015:3012],
                  prg3[3007:3004],prg3[2999:2996],prg3[2991:2988],prg3[2983:2980],prg3[2975:2972],prg3[2967:2964],prg3[2959:2956],prg3[2951:2948],
                  prg3[2943:2940],prg3[2935:2932],prg3[2927:2924],prg3[2919:2916],prg3[2911:2908],prg3[2903:2900],prg3[2895:2892],prg3[2887:2884],
                  prg3[2879:2876],prg3[2871:2868],prg3[2863:2860],prg3[2855:2852],prg3[2847:2844],prg3[2839:2836],prg3[2831:2828],prg3[2823:2820],
                  prg3[2815:2812],prg3[2807:2804],prg3[2799:2796],prg3[2791:2788],prg3[2783:2780],prg3[2775:2772],prg3[2767:2764],prg3[2759:2756],
                  prg3[2751:2748],prg3[2743:2740],prg3[2735:2732],prg3[2727:2724],prg3[2719:2716],prg3[2711:2708],prg3[2703:2700],prg3[2695:2692],
                  prg3[2687:2684],prg3[2679:2676],prg3[2671:2668],prg3[2663:2660],prg3[2655:2652],prg3[2647:2644],prg3[2639:2636],prg3[2631:2628],
                  prg3[2623:2620],prg3[2615:2612],prg3[2607:2604],prg3[2599:2596],prg3[2591:2588],prg3[2583:2580],prg3[2575:2572],prg3[2567:2564],
                  prg3[2559:2556],prg3[2551:2548],prg3[2543:2540],prg3[2535:2532],prg3[2527:2524],prg3[2519:2516],prg3[2511:2508],prg3[2503:2500],
                  prg3[2495:2492],prg3[2487:2484],prg3[2479:2476],prg3[2471:2468],prg3[2463:2460],prg3[2455:2452],prg3[2447:2444],prg3[2439:2436],
                  prg3[2431:2428],prg3[2423:2420],prg3[2415:2412],prg3[2407:2404],prg3[2399:2396],prg3[2391:2388],prg3[2383:2380],prg3[2375:2372],
                  prg3[2367:2364],prg3[2359:2356],prg3[2351:2348],prg3[2343:2340],prg3[2335:2332],prg3[2327:2324],prg3[2319:2316],prg3[2311:2308],
                  prg3[2303:2300],prg3[2295:2292],prg3[2287:2284],prg3[2279:2276],prg3[2271:2268],prg3[2263:2260],prg3[2255:2252],prg3[2247:2244],
                  prg3[2239:2236],prg3[2231:2228],prg3[2223:2220],prg3[2215:2212],prg3[2207:2204],prg3[2199:2196],prg3[2191:2188],prg3[2183:2180],
                  prg3[2175:2172],prg3[2167:2164],prg3[2159:2156],prg3[2151:2148],prg3[2143:2140],prg3[2135:2132],prg3[2127:2124],prg3[2119:2116],
                  prg3[2111:2108],prg3[2103:2100],prg3[2095:2092],prg3[2087:2084],prg3[2079:2076],prg3[2071:2068],prg3[2063:2060],prg3[2055:2052],
                  prg3[2047:2044],prg3[2039:2036],prg3[2031:2028],prg3[2023:2020],prg3[2015:2012],prg3[2007:2004],prg3[1999:1996],prg3[1991:1988],
                  prg3[1983:1980],prg3[1975:1972],prg3[1967:1964],prg3[1959:1956],prg3[1951:1948],prg3[1943:1940],prg3[1935:1932],prg3[1927:1924],
                  prg3[1919:1916],prg3[1911:1908],prg3[1903:1900],prg3[1895:1892],prg3[1887:1884],prg3[1879:1876],prg3[1871:1868],prg3[1863:1860],
                  prg3[1855:1852],prg3[1847:1844],prg3[1839:1836],prg3[1831:1828],prg3[1823:1820],prg3[1815:1812],prg3[1807:1804],prg3[1799:1796],
                  prg3[1791:1788],prg3[1783:1780],prg3[1775:1772],prg3[1767:1764],prg3[1759:1756],prg3[1751:1748],prg3[1743:1740],prg3[1735:1732],
                  prg3[1727:1724],prg3[1719:1716],prg3[1711:1708],prg3[1703:1700],prg3[1695:1692],prg3[1687:1684],prg3[1679:1676],prg3[1671:1668],
                  prg3[1663:1660],prg3[1655:1652],prg3[1647:1644],prg3[1639:1636],prg3[1631:1628],prg3[1623:1620],prg3[1615:1612],prg3[1607:1604],
                  prg3[1599:1596],prg3[1591:1588],prg3[1583:1580],prg3[1575:1572],prg3[1567:1564],prg3[1559:1556],prg3[1551:1548],prg3[1543:1540],
                  prg3[1535:1532],prg3[1527:1524],prg3[1519:1516],prg3[1511:1508],prg3[1503:1500],prg3[1495:1492],prg3[1487:1484],prg3[1479:1476],
                  prg3[1471:1468],prg3[1463:1460],prg3[1455:1452],prg3[1447:1444],prg3[1439:1436],prg3[1431:1428],prg3[1423:1420],prg3[1415:1412],
                  prg3[1407:1404],prg3[1399:1396],prg3[1391:1388],prg3[1383:1380],prg3[1375:1372],prg3[1367:1364],prg3[1359:1356],prg3[1351:1348],
                  prg3[1343:1340],prg3[1335:1332],prg3[1327:1324],prg3[1319:1316],prg3[1311:1308],prg3[1303:1300],prg3[1295:1292],prg3[1287:1284],
                  prg3[1279:1276],prg3[1271:1268],prg3[1263:1260],prg3[1255:1252],prg3[1247:1244],prg3[1239:1236],prg3[1231:1228],prg3[1223:1220],
                  prg3[1215:1212],prg3[1207:1204],prg3[1199:1196],prg3[1191:1188],prg3[1183:1180],prg3[1175:1172],prg3[1167:1164],prg3[1159:1156],
                  prg3[1151:1148],prg3[1143:1140],prg3[1135:1132],prg3[1127:1124],prg3[1119:1116],prg3[1111:1108],prg3[1103:1100],prg3[1095:1092],
                  prg3[1087:1084],prg3[1079:1076],prg3[1071:1068],prg3[1063:1060],prg3[1055:1052],prg3[1047:1044],prg3[1039:1036],prg3[1031:1028],
                  prg3[1023:1020],prg3[1015:1012],prg3[1007:1004],prg3[ 999: 996],prg3[ 991: 988],prg3[ 983: 980],prg3[ 975: 972],prg3[ 967: 964],
                  prg3[ 959: 956],prg3[ 951: 948],prg3[ 943: 940],prg3[ 935: 932],prg3[ 927: 924],prg3[ 919: 916],prg3[ 911: 908],prg3[ 903: 900],
                  prg3[ 895: 892],prg3[ 887: 884],prg3[ 879: 876],prg3[ 871: 868],prg3[ 863: 860],prg3[ 855: 852],prg3[ 847: 844],prg3[ 839: 836],
                  prg3[ 831: 828],prg3[ 823: 820],prg3[ 815: 812],prg3[ 807: 804],prg3[ 799: 796],prg3[ 791: 788],prg3[ 783: 780],prg3[ 775: 772],
                  prg3[ 767: 764],prg3[ 759: 756],prg3[ 751: 748],prg3[ 743: 740],prg3[ 735: 732],prg3[ 727: 724],prg3[ 719: 716],prg3[ 711: 708],
                  prg3[ 703: 700],prg3[ 695: 692],prg3[ 687: 684],prg3[ 679: 676],prg3[ 671: 668],prg3[ 663: 660],prg3[ 655: 652],prg3[ 647: 644],
                  prg3[ 639: 636],prg3[ 631: 628],prg3[ 623: 620],prg3[ 615: 612],prg3[ 607: 604],prg3[ 599: 596],prg3[ 591: 588],prg3[ 583: 580],
                  prg3[ 575: 572],prg3[ 567: 564],prg3[ 559: 556],prg3[ 551: 548],prg3[ 543: 540],prg3[ 535: 532],prg3[ 527: 524],prg3[ 519: 516],
                  prg3[ 511: 508],prg3[ 503: 500],prg3[ 495: 492],prg3[ 487: 484],prg3[ 479: 476],prg3[ 471: 468],prg3[ 463: 460],prg3[ 455: 452],
                  prg3[ 447: 444],prg3[ 439: 436],prg3[ 431: 428],prg3[ 423: 420],prg3[ 415: 412],prg3[ 407: 404],prg3[ 399: 396],prg3[ 391: 388],
                  prg3[ 383: 380],prg3[ 375: 372],prg3[ 367: 364],prg3[ 359: 356],prg3[ 351: 348],prg3[ 343: 340],prg3[ 335: 332],prg3[ 327: 324],
                  prg3[ 319: 316],prg3[ 311: 308],prg3[ 303: 300],prg3[ 295: 292],prg3[ 287: 284],prg3[ 279: 276],prg3[ 271: 268],prg3[ 263: 260],
                  prg3[ 255: 252],prg3[ 247: 244],prg3[ 239: 236],prg3[ 231: 228],prg3[ 223: 220],prg3[ 215: 212],prg3[ 207: 204],prg3[ 199: 196],
                  prg3[ 191: 188],prg3[ 183: 180],prg3[ 175: 172],prg3[ 167: 164],prg3[ 159: 156],prg3[ 151: 148],prg3[ 143: 140],prg3[ 135: 132],
                  prg3[ 127: 124],prg3[ 119: 116],prg3[ 111: 108],prg3[ 103: 100],prg3[  95:  92],prg3[  87:  84],prg3[  79:  76],prg3[  71:  68],
                  prg3[  63:  60],prg3[  55:  52],prg3[  47:  44],prg3[  39:  36],prg3[  31:  28],prg3[  23:  20],prg3[  15:  12],prg3[   7:   4],
                  prg2[4095:4092],prg2[4087:4084],prg2[4079:4076],prg2[4071:4068],prg2[4063:4060],prg2[4055:4052],prg2[4047:4044],prg2[4039:4036],
                  prg2[4031:4028],prg2[4023:4020],prg2[4015:4012],prg2[4007:4004],prg2[3999:3996],prg2[3991:3988],prg2[3983:3980],prg2[3975:3972],
                  prg2[3967:3964],prg2[3959:3956],prg2[3951:3948],prg2[3943:3940],prg2[3935:3932],prg2[3927:3924],prg2[3919:3916],prg2[3911:3908],
                  prg2[3903:3900],prg2[3895:3892],prg2[3887:3884],prg2[3879:3876],prg2[3871:3868],prg2[3863:3860],prg2[3855:3852],prg2[3847:3844],
                  prg2[3839:3836],prg2[3831:3828],prg2[3823:3820],prg2[3815:3812],prg2[3807:3804],prg2[3799:3796],prg2[3791:3788],prg2[3783:3780],
                  prg2[3775:3772],prg2[3767:3764],prg2[3759:3756],prg2[3751:3748],prg2[3743:3740],prg2[3735:3732],prg2[3727:3724],prg2[3719:3716],
                  prg2[3711:3708],prg2[3703:3700],prg2[3695:3692],prg2[3687:3684],prg2[3679:3676],prg2[3671:3668],prg2[3663:3660],prg2[3655:3652],
                  prg2[3647:3644],prg2[3639:3636],prg2[3631:3628],prg2[3623:3620],prg2[3615:3612],prg2[3607:3604],prg2[3599:3596],prg2[3591:3588],
                  prg2[3583:3580],prg2[3575:3572],prg2[3567:3564],prg2[3559:3556],prg2[3551:3548],prg2[3543:3540],prg2[3535:3532],prg2[3527:3524],
                  prg2[3519:3516],prg2[3511:3508],prg2[3503:3500],prg2[3495:3492],prg2[3487:3484],prg2[3479:3476],prg2[3471:3468],prg2[3463:3460],
                  prg2[3455:3452],prg2[3447:3444],prg2[3439:3436],prg2[3431:3428],prg2[3423:3420],prg2[3415:3412],prg2[3407:3404],prg2[3399:3396],
                  prg2[3391:3388],prg2[3383:3380],prg2[3375:3372],prg2[3367:3364],prg2[3359:3356],prg2[3351:3348],prg2[3343:3340],prg2[3335:3332],
                  prg2[3327:3324],prg2[3319:3316],prg2[3311:3308],prg2[3303:3300],prg2[3295:3292],prg2[3287:3284],prg2[3279:3276],prg2[3271:3268],
                  prg2[3263:3260],prg2[3255:3252],prg2[3247:3244],prg2[3239:3236],prg2[3231:3228],prg2[3223:3220],prg2[3215:3212],prg2[3207:3204],
                  prg2[3199:3196],prg2[3191:3188],prg2[3183:3180],prg2[3175:3172],prg2[3167:3164],prg2[3159:3156],prg2[3151:3148],prg2[3143:3140],
                  prg2[3135:3132],prg2[3127:3124],prg2[3119:3116],prg2[3111:3108],prg2[3103:3100],prg2[3095:3092],prg2[3087:3084],prg2[3079:3076],
                  prg2[3071:3068],prg2[3063:3060],prg2[3055:3052],prg2[3047:3044],prg2[3039:3036],prg2[3031:3028],prg2[3023:3020],prg2[3015:3012],
                  prg2[3007:3004],prg2[2999:2996],prg2[2991:2988],prg2[2983:2980],prg2[2975:2972],prg2[2967:2964],prg2[2959:2956],prg2[2951:2948],
                  prg2[2943:2940],prg2[2935:2932],prg2[2927:2924],prg2[2919:2916],prg2[2911:2908],prg2[2903:2900],prg2[2895:2892],prg2[2887:2884],
                  prg2[2879:2876],prg2[2871:2868],prg2[2863:2860],prg2[2855:2852],prg2[2847:2844],prg2[2839:2836],prg2[2831:2828],prg2[2823:2820],
                  prg2[2815:2812],prg2[2807:2804],prg2[2799:2796],prg2[2791:2788],prg2[2783:2780],prg2[2775:2772],prg2[2767:2764],prg2[2759:2756],
                  prg2[2751:2748],prg2[2743:2740],prg2[2735:2732],prg2[2727:2724],prg2[2719:2716],prg2[2711:2708],prg2[2703:2700],prg2[2695:2692],
                  prg2[2687:2684],prg2[2679:2676],prg2[2671:2668],prg2[2663:2660],prg2[2655:2652],prg2[2647:2644],prg2[2639:2636],prg2[2631:2628],
                  prg2[2623:2620],prg2[2615:2612],prg2[2607:2604],prg2[2599:2596],prg2[2591:2588],prg2[2583:2580],prg2[2575:2572],prg2[2567:2564],
                  prg2[2559:2556],prg2[2551:2548],prg2[2543:2540],prg2[2535:2532],prg2[2527:2524],prg2[2519:2516],prg2[2511:2508],prg2[2503:2500],
                  prg2[2495:2492],prg2[2487:2484],prg2[2479:2476],prg2[2471:2468],prg2[2463:2460],prg2[2455:2452],prg2[2447:2444],prg2[2439:2436],
                  prg2[2431:2428],prg2[2423:2420],prg2[2415:2412],prg2[2407:2404],prg2[2399:2396],prg2[2391:2388],prg2[2383:2380],prg2[2375:2372],
                  prg2[2367:2364],prg2[2359:2356],prg2[2351:2348],prg2[2343:2340],prg2[2335:2332],prg2[2327:2324],prg2[2319:2316],prg2[2311:2308],
                  prg2[2303:2300],prg2[2295:2292],prg2[2287:2284],prg2[2279:2276],prg2[2271:2268],prg2[2263:2260],prg2[2255:2252],prg2[2247:2244],
                  prg2[2239:2236],prg2[2231:2228],prg2[2223:2220],prg2[2215:2212],prg2[2207:2204],prg2[2199:2196],prg2[2191:2188],prg2[2183:2180],
                  prg2[2175:2172],prg2[2167:2164],prg2[2159:2156],prg2[2151:2148],prg2[2143:2140],prg2[2135:2132],prg2[2127:2124],prg2[2119:2116],
                  prg2[2111:2108],prg2[2103:2100],prg2[2095:2092],prg2[2087:2084],prg2[2079:2076],prg2[2071:2068],prg2[2063:2060],prg2[2055:2052],
                  prg2[2047:2044],prg2[2039:2036],prg2[2031:2028],prg2[2023:2020],prg2[2015:2012],prg2[2007:2004],prg2[1999:1996],prg2[1991:1988],
                  prg2[1983:1980],prg2[1975:1972],prg2[1967:1964],prg2[1959:1956],prg2[1951:1948],prg2[1943:1940],prg2[1935:1932],prg2[1927:1924],
                  prg2[1919:1916],prg2[1911:1908],prg2[1903:1900],prg2[1895:1892],prg2[1887:1884],prg2[1879:1876],prg2[1871:1868],prg2[1863:1860],
                  prg2[1855:1852],prg2[1847:1844],prg2[1839:1836],prg2[1831:1828],prg2[1823:1820],prg2[1815:1812],prg2[1807:1804],prg2[1799:1796],
                  prg2[1791:1788],prg2[1783:1780],prg2[1775:1772],prg2[1767:1764],prg2[1759:1756],prg2[1751:1748],prg2[1743:1740],prg2[1735:1732],
                  prg2[1727:1724],prg2[1719:1716],prg2[1711:1708],prg2[1703:1700],prg2[1695:1692],prg2[1687:1684],prg2[1679:1676],prg2[1671:1668],
                  prg2[1663:1660],prg2[1655:1652],prg2[1647:1644],prg2[1639:1636],prg2[1631:1628],prg2[1623:1620],prg2[1615:1612],prg2[1607:1604],
                  prg2[1599:1596],prg2[1591:1588],prg2[1583:1580],prg2[1575:1572],prg2[1567:1564],prg2[1559:1556],prg2[1551:1548],prg2[1543:1540],
                  prg2[1535:1532],prg2[1527:1524],prg2[1519:1516],prg2[1511:1508],prg2[1503:1500],prg2[1495:1492],prg2[1487:1484],prg2[1479:1476],
                  prg2[1471:1468],prg2[1463:1460],prg2[1455:1452],prg2[1447:1444],prg2[1439:1436],prg2[1431:1428],prg2[1423:1420],prg2[1415:1412],
                  prg2[1407:1404],prg2[1399:1396],prg2[1391:1388],prg2[1383:1380],prg2[1375:1372],prg2[1367:1364],prg2[1359:1356],prg2[1351:1348],
                  prg2[1343:1340],prg2[1335:1332],prg2[1327:1324],prg2[1319:1316],prg2[1311:1308],prg2[1303:1300],prg2[1295:1292],prg2[1287:1284],
                  prg2[1279:1276],prg2[1271:1268],prg2[1263:1260],prg2[1255:1252],prg2[1247:1244],prg2[1239:1236],prg2[1231:1228],prg2[1223:1220],
                  prg2[1215:1212],prg2[1207:1204],prg2[1199:1196],prg2[1191:1188],prg2[1183:1180],prg2[1175:1172],prg2[1167:1164],prg2[1159:1156],
                  prg2[1151:1148],prg2[1143:1140],prg2[1135:1132],prg2[1127:1124],prg2[1119:1116],prg2[1111:1108],prg2[1103:1100],prg2[1095:1092],
                  prg2[1087:1084],prg2[1079:1076],prg2[1071:1068],prg2[1063:1060],prg2[1055:1052],prg2[1047:1044],prg2[1039:1036],prg2[1031:1028],
                  prg2[1023:1020],prg2[1015:1012],prg2[1007:1004],prg2[ 999: 996],prg2[ 991: 988],prg2[ 983: 980],prg2[ 975: 972],prg2[ 967: 964],
                  prg2[ 959: 956],prg2[ 951: 948],prg2[ 943: 940],prg2[ 935: 932],prg2[ 927: 924],prg2[ 919: 916],prg2[ 911: 908],prg2[ 903: 900],
                  prg2[ 895: 892],prg2[ 887: 884],prg2[ 879: 876],prg2[ 871: 868],prg2[ 863: 860],prg2[ 855: 852],prg2[ 847: 844],prg2[ 839: 836],
                  prg2[ 831: 828],prg2[ 823: 820],prg2[ 815: 812],prg2[ 807: 804],prg2[ 799: 796],prg2[ 791: 788],prg2[ 783: 780],prg2[ 775: 772],
                  prg2[ 767: 764],prg2[ 759: 756],prg2[ 751: 748],prg2[ 743: 740],prg2[ 735: 732],prg2[ 727: 724],prg2[ 719: 716],prg2[ 711: 708],
                  prg2[ 703: 700],prg2[ 695: 692],prg2[ 687: 684],prg2[ 679: 676],prg2[ 671: 668],prg2[ 663: 660],prg2[ 655: 652],prg2[ 647: 644],
                  prg2[ 639: 636],prg2[ 631: 628],prg2[ 623: 620],prg2[ 615: 612],prg2[ 607: 604],prg2[ 599: 596],prg2[ 591: 588],prg2[ 583: 580],
                  prg2[ 575: 572],prg2[ 567: 564],prg2[ 559: 556],prg2[ 551: 548],prg2[ 543: 540],prg2[ 535: 532],prg2[ 527: 524],prg2[ 519: 516],
                  prg2[ 511: 508],prg2[ 503: 500],prg2[ 495: 492],prg2[ 487: 484],prg2[ 479: 476],prg2[ 471: 468],prg2[ 463: 460],prg2[ 455: 452],
                  prg2[ 447: 444],prg2[ 439: 436],prg2[ 431: 428],prg2[ 423: 420],prg2[ 415: 412],prg2[ 407: 404],prg2[ 399: 396],prg2[ 391: 388],
                  prg2[ 383: 380],prg2[ 375: 372],prg2[ 367: 364],prg2[ 359: 356],prg2[ 351: 348],prg2[ 343: 340],prg2[ 335: 332],prg2[ 327: 324],
                  prg2[ 319: 316],prg2[ 311: 308],prg2[ 303: 300],prg2[ 295: 292],prg2[ 287: 284],prg2[ 279: 276],prg2[ 271: 268],prg2[ 263: 260],
                  prg2[ 255: 252],prg2[ 247: 244],prg2[ 239: 236],prg2[ 231: 228],prg2[ 223: 220],prg2[ 215: 212],prg2[ 207: 204],prg2[ 199: 196],
                  prg2[ 191: 188],prg2[ 183: 180],prg2[ 175: 172],prg2[ 167: 164],prg2[ 159: 156],prg2[ 151: 148],prg2[ 143: 140],prg2[ 135: 132],
                  prg2[ 127: 124],prg2[ 119: 116],prg2[ 111: 108],prg2[ 103: 100],prg2[  95:  92],prg2[  87:  84],prg2[  79:  76],prg2[  71:  68],
                  prg2[  63:  60],prg2[  55:  52],prg2[  47:  44],prg2[  39:  36],prg2[  31:  28],prg2[  23:  20],prg2[  15:  12],prg2[   7:   4]};
         localparam [4095:0]
           ph0 = {prg1[4095:4092],prg1[4087:4084],prg1[4079:4076],prg1[4071:4068],prg1[4063:4060],prg1[4055:4052],prg1[4047:4044],prg1[4039:4036],
                  prg1[4031:4028],prg1[4023:4020],prg1[4015:4012],prg1[4007:4004],prg1[3999:3996],prg1[3991:3988],prg1[3983:3980],prg1[3975:3972],
                  prg1[3967:3964],prg1[3959:3956],prg1[3951:3948],prg1[3943:3940],prg1[3935:3932],prg1[3927:3924],prg1[3919:3916],prg1[3911:3908],
                  prg1[3903:3900],prg1[3895:3892],prg1[3887:3884],prg1[3879:3876],prg1[3871:3868],prg1[3863:3860],prg1[3855:3852],prg1[3847:3844],
                  prg1[3839:3836],prg1[3831:3828],prg1[3823:3820],prg1[3815:3812],prg1[3807:3804],prg1[3799:3796],prg1[3791:3788],prg1[3783:3780],
                  prg1[3775:3772],prg1[3767:3764],prg1[3759:3756],prg1[3751:3748],prg1[3743:3740],prg1[3735:3732],prg1[3727:3724],prg1[3719:3716],
                  prg1[3711:3708],prg1[3703:3700],prg1[3695:3692],prg1[3687:3684],prg1[3679:3676],prg1[3671:3668],prg1[3663:3660],prg1[3655:3652],
                  prg1[3647:3644],prg1[3639:3636],prg1[3631:3628],prg1[3623:3620],prg1[3615:3612],prg1[3607:3604],prg1[3599:3596],prg1[3591:3588],
                  prg1[3583:3580],prg1[3575:3572],prg1[3567:3564],prg1[3559:3556],prg1[3551:3548],prg1[3543:3540],prg1[3535:3532],prg1[3527:3524],
                  prg1[3519:3516],prg1[3511:3508],prg1[3503:3500],prg1[3495:3492],prg1[3487:3484],prg1[3479:3476],prg1[3471:3468],prg1[3463:3460],
                  prg1[3455:3452],prg1[3447:3444],prg1[3439:3436],prg1[3431:3428],prg1[3423:3420],prg1[3415:3412],prg1[3407:3404],prg1[3399:3396],
                  prg1[3391:3388],prg1[3383:3380],prg1[3375:3372],prg1[3367:3364],prg1[3359:3356],prg1[3351:3348],prg1[3343:3340],prg1[3335:3332],
                  prg1[3327:3324],prg1[3319:3316],prg1[3311:3308],prg1[3303:3300],prg1[3295:3292],prg1[3287:3284],prg1[3279:3276],prg1[3271:3268],
                  prg1[3263:3260],prg1[3255:3252],prg1[3247:3244],prg1[3239:3236],prg1[3231:3228],prg1[3223:3220],prg1[3215:3212],prg1[3207:3204],
                  prg1[3199:3196],prg1[3191:3188],prg1[3183:3180],prg1[3175:3172],prg1[3167:3164],prg1[3159:3156],prg1[3151:3148],prg1[3143:3140],
                  prg1[3135:3132],prg1[3127:3124],prg1[3119:3116],prg1[3111:3108],prg1[3103:3100],prg1[3095:3092],prg1[3087:3084],prg1[3079:3076],
                  prg1[3071:3068],prg1[3063:3060],prg1[3055:3052],prg1[3047:3044],prg1[3039:3036],prg1[3031:3028],prg1[3023:3020],prg1[3015:3012],
                  prg1[3007:3004],prg1[2999:2996],prg1[2991:2988],prg1[2983:2980],prg1[2975:2972],prg1[2967:2964],prg1[2959:2956],prg1[2951:2948],
                  prg1[2943:2940],prg1[2935:2932],prg1[2927:2924],prg1[2919:2916],prg1[2911:2908],prg1[2903:2900],prg1[2895:2892],prg1[2887:2884],
                  prg1[2879:2876],prg1[2871:2868],prg1[2863:2860],prg1[2855:2852],prg1[2847:2844],prg1[2839:2836],prg1[2831:2828],prg1[2823:2820],
                  prg1[2815:2812],prg1[2807:2804],prg1[2799:2796],prg1[2791:2788],prg1[2783:2780],prg1[2775:2772],prg1[2767:2764],prg1[2759:2756],
                  prg1[2751:2748],prg1[2743:2740],prg1[2735:2732],prg1[2727:2724],prg1[2719:2716],prg1[2711:2708],prg1[2703:2700],prg1[2695:2692],
                  prg1[2687:2684],prg1[2679:2676],prg1[2671:2668],prg1[2663:2660],prg1[2655:2652],prg1[2647:2644],prg1[2639:2636],prg1[2631:2628],
                  prg1[2623:2620],prg1[2615:2612],prg1[2607:2604],prg1[2599:2596],prg1[2591:2588],prg1[2583:2580],prg1[2575:2572],prg1[2567:2564],
                  prg1[2559:2556],prg1[2551:2548],prg1[2543:2540],prg1[2535:2532],prg1[2527:2524],prg1[2519:2516],prg1[2511:2508],prg1[2503:2500],
                  prg1[2495:2492],prg1[2487:2484],prg1[2479:2476],prg1[2471:2468],prg1[2463:2460],prg1[2455:2452],prg1[2447:2444],prg1[2439:2436],
                  prg1[2431:2428],prg1[2423:2420],prg1[2415:2412],prg1[2407:2404],prg1[2399:2396],prg1[2391:2388],prg1[2383:2380],prg1[2375:2372],
                  prg1[2367:2364],prg1[2359:2356],prg1[2351:2348],prg1[2343:2340],prg1[2335:2332],prg1[2327:2324],prg1[2319:2316],prg1[2311:2308],
                  prg1[2303:2300],prg1[2295:2292],prg1[2287:2284],prg1[2279:2276],prg1[2271:2268],prg1[2263:2260],prg1[2255:2252],prg1[2247:2244],
                  prg1[2239:2236],prg1[2231:2228],prg1[2223:2220],prg1[2215:2212],prg1[2207:2204],prg1[2199:2196],prg1[2191:2188],prg1[2183:2180],
                  prg1[2175:2172],prg1[2167:2164],prg1[2159:2156],prg1[2151:2148],prg1[2143:2140],prg1[2135:2132],prg1[2127:2124],prg1[2119:2116],
                  prg1[2111:2108],prg1[2103:2100],prg1[2095:2092],prg1[2087:2084],prg1[2079:2076],prg1[2071:2068],prg1[2063:2060],prg1[2055:2052],
                  prg1[2047:2044],prg1[2039:2036],prg1[2031:2028],prg1[2023:2020],prg1[2015:2012],prg1[2007:2004],prg1[1999:1996],prg1[1991:1988],
                  prg1[1983:1980],prg1[1975:1972],prg1[1967:1964],prg1[1959:1956],prg1[1951:1948],prg1[1943:1940],prg1[1935:1932],prg1[1927:1924],
                  prg1[1919:1916],prg1[1911:1908],prg1[1903:1900],prg1[1895:1892],prg1[1887:1884],prg1[1879:1876],prg1[1871:1868],prg1[1863:1860],
                  prg1[1855:1852],prg1[1847:1844],prg1[1839:1836],prg1[1831:1828],prg1[1823:1820],prg1[1815:1812],prg1[1807:1804],prg1[1799:1796],
                  prg1[1791:1788],prg1[1783:1780],prg1[1775:1772],prg1[1767:1764],prg1[1759:1756],prg1[1751:1748],prg1[1743:1740],prg1[1735:1732],
                  prg1[1727:1724],prg1[1719:1716],prg1[1711:1708],prg1[1703:1700],prg1[1695:1692],prg1[1687:1684],prg1[1679:1676],prg1[1671:1668],
                  prg1[1663:1660],prg1[1655:1652],prg1[1647:1644],prg1[1639:1636],prg1[1631:1628],prg1[1623:1620],prg1[1615:1612],prg1[1607:1604],
                  prg1[1599:1596],prg1[1591:1588],prg1[1583:1580],prg1[1575:1572],prg1[1567:1564],prg1[1559:1556],prg1[1551:1548],prg1[1543:1540],
                  prg1[1535:1532],prg1[1527:1524],prg1[1519:1516],prg1[1511:1508],prg1[1503:1500],prg1[1495:1492],prg1[1487:1484],prg1[1479:1476],
                  prg1[1471:1468],prg1[1463:1460],prg1[1455:1452],prg1[1447:1444],prg1[1439:1436],prg1[1431:1428],prg1[1423:1420],prg1[1415:1412],
                  prg1[1407:1404],prg1[1399:1396],prg1[1391:1388],prg1[1383:1380],prg1[1375:1372],prg1[1367:1364],prg1[1359:1356],prg1[1351:1348],
                  prg1[1343:1340],prg1[1335:1332],prg1[1327:1324],prg1[1319:1316],prg1[1311:1308],prg1[1303:1300],prg1[1295:1292],prg1[1287:1284],
                  prg1[1279:1276],prg1[1271:1268],prg1[1263:1260],prg1[1255:1252],prg1[1247:1244],prg1[1239:1236],prg1[1231:1228],prg1[1223:1220],
                  prg1[1215:1212],prg1[1207:1204],prg1[1199:1196],prg1[1191:1188],prg1[1183:1180],prg1[1175:1172],prg1[1167:1164],prg1[1159:1156],
                  prg1[1151:1148],prg1[1143:1140],prg1[1135:1132],prg1[1127:1124],prg1[1119:1116],prg1[1111:1108],prg1[1103:1100],prg1[1095:1092],
                  prg1[1087:1084],prg1[1079:1076],prg1[1071:1068],prg1[1063:1060],prg1[1055:1052],prg1[1047:1044],prg1[1039:1036],prg1[1031:1028],
                  prg1[1023:1020],prg1[1015:1012],prg1[1007:1004],prg1[ 999: 996],prg1[ 991: 988],prg1[ 983: 980],prg1[ 975: 972],prg1[ 967: 964],
                  prg1[ 959: 956],prg1[ 951: 948],prg1[ 943: 940],prg1[ 935: 932],prg1[ 927: 924],prg1[ 919: 916],prg1[ 911: 908],prg1[ 903: 900],
                  prg1[ 895: 892],prg1[ 887: 884],prg1[ 879: 876],prg1[ 871: 868],prg1[ 863: 860],prg1[ 855: 852],prg1[ 847: 844],prg1[ 839: 836],
                  prg1[ 831: 828],prg1[ 823: 820],prg1[ 815: 812],prg1[ 807: 804],prg1[ 799: 796],prg1[ 791: 788],prg1[ 783: 780],prg1[ 775: 772],
                  prg1[ 767: 764],prg1[ 759: 756],prg1[ 751: 748],prg1[ 743: 740],prg1[ 735: 732],prg1[ 727: 724],prg1[ 719: 716],prg1[ 711: 708],
                  prg1[ 703: 700],prg1[ 695: 692],prg1[ 687: 684],prg1[ 679: 676],prg1[ 671: 668],prg1[ 663: 660],prg1[ 655: 652],prg1[ 647: 644],
                  prg1[ 639: 636],prg1[ 631: 628],prg1[ 623: 620],prg1[ 615: 612],prg1[ 607: 604],prg1[ 599: 596],prg1[ 591: 588],prg1[ 583: 580],
                  prg1[ 575: 572],prg1[ 567: 564],prg1[ 559: 556],prg1[ 551: 548],prg1[ 543: 540],prg1[ 535: 532],prg1[ 527: 524],prg1[ 519: 516],
                  prg1[ 511: 508],prg1[ 503: 500],prg1[ 495: 492],prg1[ 487: 484],prg1[ 479: 476],prg1[ 471: 468],prg1[ 463: 460],prg1[ 455: 452],
                  prg1[ 447: 444],prg1[ 439: 436],prg1[ 431: 428],prg1[ 423: 420],prg1[ 415: 412],prg1[ 407: 404],prg1[ 399: 396],prg1[ 391: 388],
                  prg1[ 383: 380],prg1[ 375: 372],prg1[ 367: 364],prg1[ 359: 356],prg1[ 351: 348],prg1[ 343: 340],prg1[ 335: 332],prg1[ 327: 324],
                  prg1[ 319: 316],prg1[ 311: 308],prg1[ 303: 300],prg1[ 295: 292],prg1[ 287: 284],prg1[ 279: 276],prg1[ 271: 268],prg1[ 263: 260],
                  prg1[ 255: 252],prg1[ 247: 244],prg1[ 239: 236],prg1[ 231: 228],prg1[ 223: 220],prg1[ 215: 212],prg1[ 207: 204],prg1[ 199: 196],
                  prg1[ 191: 188],prg1[ 183: 180],prg1[ 175: 172],prg1[ 167: 164],prg1[ 159: 156],prg1[ 151: 148],prg1[ 143: 140],prg1[ 135: 132],
                  prg1[ 127: 124],prg1[ 119: 116],prg1[ 111: 108],prg1[ 103: 100],prg1[  95:  92],prg1[  87:  84],prg1[  79:  76],prg1[  71:  68],
                  prg1[  63:  60],prg1[  55:  52],prg1[  47:  44],prg1[  39:  36],prg1[  31:  28],prg1[  23:  20],prg1[  15:  12],prg1[   7:   4],
                  prg0[4095:4092],prg0[4087:4084],prg0[4079:4076],prg0[4071:4068],prg0[4063:4060],prg0[4055:4052],prg0[4047:4044],prg0[4039:4036],
                  prg0[4031:4028],prg0[4023:4020],prg0[4015:4012],prg0[4007:4004],prg0[3999:3996],prg0[3991:3988],prg0[3983:3980],prg0[3975:3972],
                  prg0[3967:3964],prg0[3959:3956],prg0[3951:3948],prg0[3943:3940],prg0[3935:3932],prg0[3927:3924],prg0[3919:3916],prg0[3911:3908],
                  prg0[3903:3900],prg0[3895:3892],prg0[3887:3884],prg0[3879:3876],prg0[3871:3868],prg0[3863:3860],prg0[3855:3852],prg0[3847:3844],
                  prg0[3839:3836],prg0[3831:3828],prg0[3823:3820],prg0[3815:3812],prg0[3807:3804],prg0[3799:3796],prg0[3791:3788],prg0[3783:3780],
                  prg0[3775:3772],prg0[3767:3764],prg0[3759:3756],prg0[3751:3748],prg0[3743:3740],prg0[3735:3732],prg0[3727:3724],prg0[3719:3716],
                  prg0[3711:3708],prg0[3703:3700],prg0[3695:3692],prg0[3687:3684],prg0[3679:3676],prg0[3671:3668],prg0[3663:3660],prg0[3655:3652],
                  prg0[3647:3644],prg0[3639:3636],prg0[3631:3628],prg0[3623:3620],prg0[3615:3612],prg0[3607:3604],prg0[3599:3596],prg0[3591:3588],
                  prg0[3583:3580],prg0[3575:3572],prg0[3567:3564],prg0[3559:3556],prg0[3551:3548],prg0[3543:3540],prg0[3535:3532],prg0[3527:3524],
                  prg0[3519:3516],prg0[3511:3508],prg0[3503:3500],prg0[3495:3492],prg0[3487:3484],prg0[3479:3476],prg0[3471:3468],prg0[3463:3460],
                  prg0[3455:3452],prg0[3447:3444],prg0[3439:3436],prg0[3431:3428],prg0[3423:3420],prg0[3415:3412],prg0[3407:3404],prg0[3399:3396],
                  prg0[3391:3388],prg0[3383:3380],prg0[3375:3372],prg0[3367:3364],prg0[3359:3356],prg0[3351:3348],prg0[3343:3340],prg0[3335:3332],
                  prg0[3327:3324],prg0[3319:3316],prg0[3311:3308],prg0[3303:3300],prg0[3295:3292],prg0[3287:3284],prg0[3279:3276],prg0[3271:3268],
                  prg0[3263:3260],prg0[3255:3252],prg0[3247:3244],prg0[3239:3236],prg0[3231:3228],prg0[3223:3220],prg0[3215:3212],prg0[3207:3204],
                  prg0[3199:3196],prg0[3191:3188],prg0[3183:3180],prg0[3175:3172],prg0[3167:3164],prg0[3159:3156],prg0[3151:3148],prg0[3143:3140],
                  prg0[3135:3132],prg0[3127:3124],prg0[3119:3116],prg0[3111:3108],prg0[3103:3100],prg0[3095:3092],prg0[3087:3084],prg0[3079:3076],
                  prg0[3071:3068],prg0[3063:3060],prg0[3055:3052],prg0[3047:3044],prg0[3039:3036],prg0[3031:3028],prg0[3023:3020],prg0[3015:3012],
                  prg0[3007:3004],prg0[2999:2996],prg0[2991:2988],prg0[2983:2980],prg0[2975:2972],prg0[2967:2964],prg0[2959:2956],prg0[2951:2948],
                  prg0[2943:2940],prg0[2935:2932],prg0[2927:2924],prg0[2919:2916],prg0[2911:2908],prg0[2903:2900],prg0[2895:2892],prg0[2887:2884],
                  prg0[2879:2876],prg0[2871:2868],prg0[2863:2860],prg0[2855:2852],prg0[2847:2844],prg0[2839:2836],prg0[2831:2828],prg0[2823:2820],
                  prg0[2815:2812],prg0[2807:2804],prg0[2799:2796],prg0[2791:2788],prg0[2783:2780],prg0[2775:2772],prg0[2767:2764],prg0[2759:2756],
                  prg0[2751:2748],prg0[2743:2740],prg0[2735:2732],prg0[2727:2724],prg0[2719:2716],prg0[2711:2708],prg0[2703:2700],prg0[2695:2692],
                  prg0[2687:2684],prg0[2679:2676],prg0[2671:2668],prg0[2663:2660],prg0[2655:2652],prg0[2647:2644],prg0[2639:2636],prg0[2631:2628],
                  prg0[2623:2620],prg0[2615:2612],prg0[2607:2604],prg0[2599:2596],prg0[2591:2588],prg0[2583:2580],prg0[2575:2572],prg0[2567:2564],
                  prg0[2559:2556],prg0[2551:2548],prg0[2543:2540],prg0[2535:2532],prg0[2527:2524],prg0[2519:2516],prg0[2511:2508],prg0[2503:2500],
                  prg0[2495:2492],prg0[2487:2484],prg0[2479:2476],prg0[2471:2468],prg0[2463:2460],prg0[2455:2452],prg0[2447:2444],prg0[2439:2436],
                  prg0[2431:2428],prg0[2423:2420],prg0[2415:2412],prg0[2407:2404],prg0[2399:2396],prg0[2391:2388],prg0[2383:2380],prg0[2375:2372],
                  prg0[2367:2364],prg0[2359:2356],prg0[2351:2348],prg0[2343:2340],prg0[2335:2332],prg0[2327:2324],prg0[2319:2316],prg0[2311:2308],
                  prg0[2303:2300],prg0[2295:2292],prg0[2287:2284],prg0[2279:2276],prg0[2271:2268],prg0[2263:2260],prg0[2255:2252],prg0[2247:2244],
                  prg0[2239:2236],prg0[2231:2228],prg0[2223:2220],prg0[2215:2212],prg0[2207:2204],prg0[2199:2196],prg0[2191:2188],prg0[2183:2180],
                  prg0[2175:2172],prg0[2167:2164],prg0[2159:2156],prg0[2151:2148],prg0[2143:2140],prg0[2135:2132],prg0[2127:2124],prg0[2119:2116],
                  prg0[2111:2108],prg0[2103:2100],prg0[2095:2092],prg0[2087:2084],prg0[2079:2076],prg0[2071:2068],prg0[2063:2060],prg0[2055:2052],
                  prg0[2047:2044],prg0[2039:2036],prg0[2031:2028],prg0[2023:2020],prg0[2015:2012],prg0[2007:2004],prg0[1999:1996],prg0[1991:1988],
                  prg0[1983:1980],prg0[1975:1972],prg0[1967:1964],prg0[1959:1956],prg0[1951:1948],prg0[1943:1940],prg0[1935:1932],prg0[1927:1924],
                  prg0[1919:1916],prg0[1911:1908],prg0[1903:1900],prg0[1895:1892],prg0[1887:1884],prg0[1879:1876],prg0[1871:1868],prg0[1863:1860],
                  prg0[1855:1852],prg0[1847:1844],prg0[1839:1836],prg0[1831:1828],prg0[1823:1820],prg0[1815:1812],prg0[1807:1804],prg0[1799:1796],
                  prg0[1791:1788],prg0[1783:1780],prg0[1775:1772],prg0[1767:1764],prg0[1759:1756],prg0[1751:1748],prg0[1743:1740],prg0[1735:1732],
                  prg0[1727:1724],prg0[1719:1716],prg0[1711:1708],prg0[1703:1700],prg0[1695:1692],prg0[1687:1684],prg0[1679:1676],prg0[1671:1668],
                  prg0[1663:1660],prg0[1655:1652],prg0[1647:1644],prg0[1639:1636],prg0[1631:1628],prg0[1623:1620],prg0[1615:1612],prg0[1607:1604],
                  prg0[1599:1596],prg0[1591:1588],prg0[1583:1580],prg0[1575:1572],prg0[1567:1564],prg0[1559:1556],prg0[1551:1548],prg0[1543:1540],
                  prg0[1535:1532],prg0[1527:1524],prg0[1519:1516],prg0[1511:1508],prg0[1503:1500],prg0[1495:1492],prg0[1487:1484],prg0[1479:1476],
                  prg0[1471:1468],prg0[1463:1460],prg0[1455:1452],prg0[1447:1444],prg0[1439:1436],prg0[1431:1428],prg0[1423:1420],prg0[1415:1412],
                  prg0[1407:1404],prg0[1399:1396],prg0[1391:1388],prg0[1383:1380],prg0[1375:1372],prg0[1367:1364],prg0[1359:1356],prg0[1351:1348],
                  prg0[1343:1340],prg0[1335:1332],prg0[1327:1324],prg0[1319:1316],prg0[1311:1308],prg0[1303:1300],prg0[1295:1292],prg0[1287:1284],
                  prg0[1279:1276],prg0[1271:1268],prg0[1263:1260],prg0[1255:1252],prg0[1247:1244],prg0[1239:1236],prg0[1231:1228],prg0[1223:1220],
                  prg0[1215:1212],prg0[1207:1204],prg0[1199:1196],prg0[1191:1188],prg0[1183:1180],prg0[1175:1172],prg0[1167:1164],prg0[1159:1156],
                  prg0[1151:1148],prg0[1143:1140],prg0[1135:1132],prg0[1127:1124],prg0[1119:1116],prg0[1111:1108],prg0[1103:1100],prg0[1095:1092],
                  prg0[1087:1084],prg0[1079:1076],prg0[1071:1068],prg0[1063:1060],prg0[1055:1052],prg0[1047:1044],prg0[1039:1036],prg0[1031:1028],
                  prg0[1023:1020],prg0[1015:1012],prg0[1007:1004],prg0[ 999: 996],prg0[ 991: 988],prg0[ 983: 980],prg0[ 975: 972],prg0[ 967: 964],
                  prg0[ 959: 956],prg0[ 951: 948],prg0[ 943: 940],prg0[ 935: 932],prg0[ 927: 924],prg0[ 919: 916],prg0[ 911: 908],prg0[ 903: 900],
                  prg0[ 895: 892],prg0[ 887: 884],prg0[ 879: 876],prg0[ 871: 868],prg0[ 863: 860],prg0[ 855: 852],prg0[ 847: 844],prg0[ 839: 836],
                  prg0[ 831: 828],prg0[ 823: 820],prg0[ 815: 812],prg0[ 807: 804],prg0[ 799: 796],prg0[ 791: 788],prg0[ 783: 780],prg0[ 775: 772],
                  prg0[ 767: 764],prg0[ 759: 756],prg0[ 751: 748],prg0[ 743: 740],prg0[ 735: 732],prg0[ 727: 724],prg0[ 719: 716],prg0[ 711: 708],
                  prg0[ 703: 700],prg0[ 695: 692],prg0[ 687: 684],prg0[ 679: 676],prg0[ 671: 668],prg0[ 663: 660],prg0[ 655: 652],prg0[ 647: 644],
                  prg0[ 639: 636],prg0[ 631: 628],prg0[ 623: 620],prg0[ 615: 612],prg0[ 607: 604],prg0[ 599: 596],prg0[ 591: 588],prg0[ 583: 580],
                  prg0[ 575: 572],prg0[ 567: 564],prg0[ 559: 556],prg0[ 551: 548],prg0[ 543: 540],prg0[ 535: 532],prg0[ 527: 524],prg0[ 519: 516],
                  prg0[ 511: 508],prg0[ 503: 500],prg0[ 495: 492],prg0[ 487: 484],prg0[ 479: 476],prg0[ 471: 468],prg0[ 463: 460],prg0[ 455: 452],
                  prg0[ 447: 444],prg0[ 439: 436],prg0[ 431: 428],prg0[ 423: 420],prg0[ 415: 412],prg0[ 407: 404],prg0[ 399: 396],prg0[ 391: 388],
                  prg0[ 383: 380],prg0[ 375: 372],prg0[ 367: 364],prg0[ 359: 356],prg0[ 351: 348],prg0[ 343: 340],prg0[ 335: 332],prg0[ 327: 324],
                  prg0[ 319: 316],prg0[ 311: 308],prg0[ 303: 300],prg0[ 295: 292],prg0[ 287: 284],prg0[ 279: 276],prg0[ 271: 268],prg0[ 263: 260],
                  prg0[ 255: 252],prg0[ 247: 244],prg0[ 239: 236],prg0[ 231: 228],prg0[ 223: 220],prg0[ 215: 212],prg0[ 207: 204],prg0[ 199: 196],
                  prg0[ 191: 188],prg0[ 183: 180],prg0[ 175: 172],prg0[ 167: 164],prg0[ 159: 156],prg0[ 151: 148],prg0[ 143: 140],prg0[ 135: 132],
                  prg0[ 127: 124],prg0[ 119: 116],prg0[ 111: 108],prg0[ 103: 100],prg0[  95:  92],prg0[  87:  84],prg0[  79:  76],prg0[  71:  68],
                  prg0[  63:  60],prg0[  55:  52],prg0[  47:  44],prg0[  39:  36],prg0[  31:  28],prg0[  23:  20],prg0[  15:  12],prg0[   7:   4]};

         m_ebr_w4 #(.EBRADRWIDTH(EBRADRWIDTH),
                    .prg0(pb0), .prg1(pb1))
         ebrb 
           (/*AUTOINST*/
            // Outputs
            .DAT_O                      (DAT_O[3:0]),
            // Inputs
            .B                          (B[3:0]),
            .Rai                        (Rai[EBRADRWIDTH-1:0]),
            .Wai                        (Wai[EBRADRWIDTH-1:0]),
            .clk                        (clk),
            .we                         (we));
   
         m_ebr_w4 #(.EBRADRWIDTH(EBRADRWIDTH),
                    .prg0(ph0), .prg1(ph1))
         ebrh 
           (// Outputs
            .DAT_O                      (DAT_O[7:4]),
            // Inputs
            .B                          (B[7:4]),
            /*AUTOINST*/
            // Inputs
            .Rai                        (Rai[EBRADRWIDTH-1:0]),
            .Wai                        (Wai[EBRADRWIDTH-1:0]),
            .clk                        (clk),
            .we                         (we));
   
      end
   endgenerate
endmodule


// Local Variables:
// verilog-library-directories:("." "sb_sim_rtl" )
// verilog-library-extensions:(".v" )
// End:
