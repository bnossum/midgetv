-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Oct 12 2020 16:05:25

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    TX : out std_logic;
    RX : in std_logic;
    LED4 : out std_logic;
    LED3 : out std_logic;
    LED2 : out std_logic;
    LED1 : out std_logic;
    CLK : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__15400\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \VCCG0\ : std_logic;
signal \inst_midgetv_core.Wai_8\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.n28\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.n5610\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_0\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_1\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_2\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_3\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_4\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_5\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_6\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_7\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_6\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_3\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_2\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_4\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa07h\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \inst_midgetv_core.inst_alu_carryin.genblk1_genblk1_prealucyin\ : std_logic;
signal \inst_midgetv_core.alu_carryin\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_1\ : std_logic;
signal \inst_midgetv_core.QQ_2\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_2\ : std_logic;
signal \inst_midgetv_core.QQ_3\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_3\ : std_logic;
signal \inst_midgetv_core.QQ_4\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_4\ : std_logic;
signal \GNDG0\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_5\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_5_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \inst_midgetv_core.QQ_6\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_6\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_7\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_8\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_9\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_10\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_11\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_12\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_13\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_14\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_15\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_16\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_17\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_18\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_19\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_20\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_21\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_22\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_23\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_24\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_25\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_26\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_27\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_28\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_29\ : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_30\ : std_logic;
signal \inst_midgetv_core.s_alu_2\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.alucy_31\ : std_logic;
signal \inst_midgetv_core.alu_carryout\ : std_logic;
signal \inst_midgetv_core.inst_condcode.n2\ : std_logic;
signal \inst_midgetv_core.alu_carryout_THRU_CO\ : std_logic;
signal \inst_midgetv_core.inst_condcode.n6\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.n5608\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.n5609\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_0\ : std_logic;
signal \inst_midgetv_core.QQ_0\ : std_logic;
signal \inst_midgetv_core.s_cyclecnt_1\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_1\ : std_logic;
signal \inst_midgetv_core.QQ_1\ : std_logic;
signal \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_5\ : std_logic;
signal \inst_midgetv_core.QQ_5\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy1\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy2\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy3\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm4a\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy4\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy5\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy6\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy7\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy8\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy9\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy10\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm11b\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm11a\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy11\ : std_logic;
signal \inst_midgetv_core.B_12\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy12\ : std_logic;
signal \inst_midgetv_core.B_13\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy13\ : std_logic;
signal \inst_midgetv_core.B_14\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy14\ : std_logic;
signal \inst_midgetv_core.B_15\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy15\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy16\ : std_logic;
signal \inst_midgetv_core.B_16\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \inst_midgetv_core.B_17\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy17\ : std_logic;
signal \inst_midgetv_core.B_18\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy18\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa13b\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa31\ : std_logic;
signal \inst_midgetv_core.B_19\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy19\ : std_logic;
signal \inst_midgetv_core.B_20\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy20\ : std_logic;
signal \inst_midgetv_core.B_21\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy21\ : std_logic;
signal \inst_midgetv_core.B_22\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy22\ : std_logic;
signal \inst_midgetv_core.B_23\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy23\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy24\ : std_logic;
signal \inst_midgetv_core.B_24\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \inst_midgetv_core.B_25\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy25\ : std_logic;
signal \inst_midgetv_core.B_26\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy26\ : std_logic;
signal \inst_midgetv_core.B_27\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy27\ : std_logic;
signal \inst_midgetv_core.B_28\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy28\ : std_logic;
signal \inst_midgetv_core.B_29\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy29\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy30\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa13\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa10\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy31\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy32\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \inst_midgetv_core.DAT_O_21\ : std_logic;
signal \inst_midgetv_core.Di_21_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_21\ : std_logic;
signal \inst_midgetv_core.DAT_O_22\ : std_logic;
signal \inst_midgetv_core.ADR_O_22\ : std_logic;
signal \inst_midgetv_core.Di_22_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_22\ : std_logic;
signal \inst_midgetv_core.DAT_O_23\ : std_logic;
signal \inst_midgetv_core.ADR_O_23\ : std_logic;
signal \inst_midgetv_core.Di_23_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_23\ : std_logic;
signal \inst_midgetv_core.DAT_O_24\ : std_logic;
signal \inst_midgetv_core.ADR_O_24\ : std_logic;
signal \inst_midgetv_core.Di_24_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_24\ : std_logic;
signal \inst_midgetv_core.Wai_7\ : std_logic;
signal \inst_midgetv_core.mostofminx0\ : std_logic;
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.instr0100\ : std_logic;
signal \inst_midgetv_core.rinx_4\ : std_logic;
signal \inst_midgetv_core.minx_4\ : std_logic;
signal \inst_midgetv_core.rinx_2\ : std_logic;
signal \inst_midgetv_core.minx_2\ : std_logic;
signal \inst_midgetv_core.sa43\ : std_logic;
signal \inst_midgetv_core.inst_progressctrl.n2764\ : std_logic;
signal \inst_midgetv_core.inst_progressctrl.ctrlreg_we_N_84\ : std_logic;
signal \inst_midgetv_core.sa14\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_nsa14_or_nCORERUNNING\ : std_logic;
signal \DAT_O_0\ : std_logic;
signal \inst_midgetv_core.INSTR_0\ : std_logic;
signal \inst_midgetv_core.ADR_O_0\ : std_logic;
signal \inst_midgetv_core.Di_0_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_0\ : std_logic;
signal \DAT_O_1\ : std_logic;
signal \inst_midgetv_core.INSTR_1\ : std_logic;
signal \inst_midgetv_core.Di_1_cascade_\ : std_logic;
signal \inst_midgetv_core.ADR_O_1\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_1\ : std_logic;
signal \inst_midgetv_core.Di_2_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_2\ : std_logic;
signal \DAT_O_3\ : std_logic;
signal \inst_midgetv_core.Di_3_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_3\ : std_logic;
signal \inst_midgetv_core.DAT_O_4\ : std_logic;
signal \inst_midgetv_core.Di_4_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_4\ : std_logic;
signal \inst_midgetv_core.DAT_O_5\ : std_logic;
signal \inst_midgetv_core.Di_5_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_5\ : std_logic;
signal \inst_midgetv_core.DAT_O_6\ : std_logic;
signal \inst_midgetv_core.Di_6_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_6\ : std_logic;
signal \inst_midgetv_core.DAT_O_8\ : std_logic;
signal \inst_midgetv_core.Di_8_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_8\ : std_logic;
signal \inst_midgetv_core.DAT_O_10\ : std_logic;
signal \inst_midgetv_core.Di_10_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_10\ : std_logic;
signal \inst_midgetv_core.DAT_O_11\ : std_logic;
signal \inst_midgetv_core.Di_11_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_11\ : std_logic;
signal \inst_midgetv_core.ADR_O_10\ : std_logic;
signal \inst_midgetv_core.DAT_O_9\ : std_logic;
signal \inst_midgetv_core.Di_9_cascade_\ : std_logic;
signal \inst_midgetv_core.ADR_O_9\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_9\ : std_logic;
signal \inst_midgetv_core.DAT_O_12\ : std_logic;
signal \inst_midgetv_core.ADR_O_12\ : std_logic;
signal \inst_midgetv_core.Di_12_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_12\ : std_logic;
signal \inst_midgetv_core.DAT_O_29\ : std_logic;
signal \inst_midgetv_core.Di_29_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_29\ : std_logic;
signal \inst_midgetv_core.DAT_O_30\ : std_logic;
signal \inst_midgetv_core.ADR_O_30\ : std_logic;
signal \inst_midgetv_core.Di_30_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_30\ : std_logic;
signal \inst_midgetv_core.sra_msb\ : std_logic;
signal \inst_midgetv_core.ADR_O_31\ : std_logic;
signal \inst_midgetv_core.Di_31_cascade_\ : std_logic;
signal \inst_midgetv_core.A31\ : std_logic;
signal \inst_midgetv_core.DAT_O_7\ : std_logic;
signal \inst_midgetv_core.Di_7_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_7\ : std_logic;
signal \inst_midgetv_core.DAT_O_17\ : std_logic;
signal \inst_midgetv_core.Di_17_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_17\ : std_logic;
signal \inst_midgetv_core.DAT_O_18\ : std_logic;
signal \inst_midgetv_core.ADR_O_18\ : std_logic;
signal \inst_midgetv_core.Di_18_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_18\ : std_logic;
signal \inst_midgetv_core.DAT_O_19\ : std_logic;
signal \inst_midgetv_core.ADR_O_19\ : std_logic;
signal \inst_midgetv_core.Di_19_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_19\ : std_logic;
signal \inst_midgetv_core.DAT_O_20\ : std_logic;
signal \inst_midgetv_core.ADR_O_21\ : std_logic;
signal \inst_midgetv_core.ADR_O_20\ : std_logic;
signal \inst_midgetv_core.Di_20_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_20\ : std_logic;
signal \inst_midgetv_core.DAT_O_25\ : std_logic;
signal \inst_midgetv_core.Di_25_cascade_\ : std_logic;
signal \inst_midgetv_core.ADR_O_25\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_25\ : std_logic;
signal \inst_midgetv_core.DAT_O_26\ : std_logic;
signal \inst_midgetv_core.ADR_O_26\ : std_logic;
signal \inst_midgetv_core.Di_26_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_26\ : std_logic;
signal \inst_midgetv_core.DAT_O_27\ : std_logic;
signal \inst_midgetv_core.ADR_O_27\ : std_logic;
signal \inst_midgetv_core.Di_27_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_27\ : std_logic;
signal \inst_midgetv_core.ADR_O_29\ : std_logic;
signal \inst_midgetv_core.DAT_O_28\ : std_logic;
signal \inst_midgetv_core.ADR_O_28\ : std_logic;
signal \inst_midgetv_core.Di_28_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_28\ : std_logic;
signal \inst_midgetv_core.rinx_1\ : std_logic;
signal \inst_midgetv_core.minx_1\ : std_logic;
signal \inst_midgetv_core.rinx_5\ : std_logic;
signal \inst_midgetv_core.minx_5\ : std_logic;
signal \inst_midgetv_core.rinx_7\ : std_logic;
signal \inst_midgetv_core.minx_7\ : std_logic;
signal \inst_midgetv_core.rinx_3\ : std_logic;
signal \inst_midgetv_core.minx_3\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.usedinx_or_RST_I_notcorerunning\ : std_logic;
signal \inst_midgetv_core.rinx_6\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.illegal\ : std_logic;
signal \inst_midgetv_core.minx_6\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.n15\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09h\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.n5603\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.n17\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.dinx_1_N_145_0\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.n5613\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk2_illegal_a\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.n6\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.n2\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk1_checkfunct7_N_286\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.n5605\ : std_logic;
signal \inst_midgetv_core.INSTR_3\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.n8\ : std_logic;
signal \inst_midgetv_core.FUNC7_2\ : std_logic;
signal \inst_midgetv_core.FUNC7_4\ : std_logic;
signal \inst_midgetv_core.FUNC7_5\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.n497\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.n11\ : std_logic;
signal \inst_midgetv_core.INSTR_5\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.n2575\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk1_checkfunct7_N_281\ : std_logic;
signal \inst_midgetv_core.raluF\ : std_logic;
signal \inst_midgetv_core.is_brcond\ : std_logic;
signal \inst_midgetv_core.rzcy32\ : std_logic;
signal \inst_midgetv_core.INSTR_12\ : std_logic;
signal \inst_midgetv_core.inst_condcode.n5618\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk1_illegal_rs1_rd_N_300\ : std_logic;
signal \uart_ACK_O\ : std_logic;
signal \rDee_8\ : std_logic;
signal \inst_midgetv_core.FUNC7_6\ : std_logic;
signal \inst_midgetv_core.FUNC7_1\ : std_logic;
signal \inst_midgetv_core.FUNC7_3\ : std_logic;
signal \inst_midgetv_core.FUNC7_0\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.n12\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.n17\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.inst_illegalop.n16\ : std_logic;
signal \inst_midgetv_core.DAT_O_13\ : std_logic;
signal \inst_midgetv_core.INSTR_13\ : std_logic;
signal \inst_midgetv_core.Di_13_cascade_\ : std_logic;
signal \inst_midgetv_core.ADR_O_13\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_13\ : std_logic;
signal \inst_midgetv_core.DAT_O_14\ : std_logic;
signal \inst_midgetv_core.INSTR_14\ : std_logic;
signal \inst_midgetv_core.ADR_O_14\ : std_logic;
signal \inst_midgetv_core.Di_14_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_14\ : std_logic;
signal \inst_midgetv_core.DAT_O_15\ : std_logic;
signal \inst_midgetv_core.ADR_O_15\ : std_logic;
signal \inst_midgetv_core.Di_15_cascade_\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_15\ : std_logic;
signal \inst_midgetv_core.ADR_O_17\ : std_logic;
signal \inst_midgetv_core.DAT_O_16\ : std_logic;
signal \inst_midgetv_core.inst_mimux.genblk1_sa00mod\ : std_logic;
signal \inst_midgetv_core.ADR_O_16\ : std_logic;
signal \inst_midgetv_core.s_alu_1\ : std_logic;
signal \inst_midgetv_core.Di_16_cascade_\ : std_logic;
signal \inst_midgetv_core.s_alu_0\ : std_logic;
signal \inst_midgetv_core.inst_alu.genblk1_inst.A_16\ : std_logic;
signal \inst_midgetv_core.B_30\ : std_logic;
signal \inst_midgetv_core.sa29\ : std_logic;
signal \inst_midgetv_core.is_valid_instrhigh\ : std_logic;
signal \inst_midgetv_core.progress_ucode\ : std_logic;
signal \inst_midgetv_core.rinx_0\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.n5624\ : std_logic;
signal \inst_midgetv_core.sa33\ : std_logic;
signal \inst_midgetv_core.inst_progressctrl.n4\ : std_logic;
signal \inst_midgetv_core.enaQ\ : std_logic;
signal \inst_midgetv_core.sa00\ : std_logic;
signal \inst_midgetv_core.Wai_0\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \inst_midgetv_core.Wai_1\ : std_logic;
signal \inst_midgetv_core.inst_wai.genblk1_waicy0\ : std_logic;
signal \inst_midgetv_core.ADR_O_4\ : std_logic;
signal \inst_midgetv_core.Wai_2\ : std_logic;
signal \inst_midgetv_core.inst_wai.genblk1_waicy1\ : std_logic;
signal \inst_midgetv_core.ADR_O_5\ : std_logic;
signal \inst_midgetv_core.Wai_3\ : std_logic;
signal \inst_midgetv_core.inst_wai.genblk1_waicy2\ : std_logic;
signal \inst_midgetv_core.INSTR_11\ : std_logic;
signal \inst_midgetv_core.ADR_O_6\ : std_logic;
signal \inst_midgetv_core.Wai_4\ : std_logic;
signal \inst_midgetv_core.inst_wai.genblk1_waicy3\ : std_logic;
signal \inst_midgetv_core.ADR_O_7\ : std_logic;
signal \inst_midgetv_core.inst_wai.genblk1_waicy4\ : std_logic;
signal \inst_midgetv_core.Wai_5\ : std_logic;
signal \inst_midgetv_core.inst_wai.genblk1_preWai0\ : std_logic;
signal \inst_midgetv_core.INSTR_7\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm0a\ : std_logic;
signal \inst_midgetv_core.INSTR_9\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm2a\ : std_logic;
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.we\ : std_logic;
signal \inst_midgetv_core.INSTR_6\ : std_logic;
signal \inst_midgetv_core.INSTR_2\ : std_logic;
signal \inst_midgetv_core.s_cyclecnt_0\ : std_logic;
signal \inst_midgetv_core.INSTR_4\ : std_logic;
signal \inst_midgetv_core.INSTR_8\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm1a\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa07\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa08\ : std_logic;
signal \inst_midgetv_core.INSTR_10\ : std_logic;
signal \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm3a\ : std_logic;
signal \inst_midgetv_core.bmask_0\ : std_logic;
signal \inst_midgetv_core.rlastshift\ : std_logic;
signal \inst_midgetv_core.sa41\ : std_logic;
signal corerunning : std_logic;
signal \inst_midgetv_core.inst_progressctrl.blka_cmb_bsel_3_cascade_\ : std_logic;
signal \meta_usartRX\ : std_logic;
signal \DAT_O_2\ : std_logic;
signal \LED3_c\ : std_logic;
signal \inst_midgetv_core.ADR_O_11\ : std_logic;
signal \inst_midgetv_core.Wai_9\ : std_logic;
signal \SEL_O_3\ : std_logic;
signal \DAT_O_31\ : std_logic;
signal bluesource_is_uart : std_logic;
signal \i_LEDs.n2766\ : std_logic;
signal \i_BBUART.usartTX_N_2\ : std_logic;
signal \WE_O\ : std_logic;
signal \ADR_O_2\ : std_logic;
signal \LED1_N_4\ : std_logic;
signal \inst_midgetv_core.inst_progressctrl.n4_adj_311\ : std_logic;
signal n2345 : std_logic;
signal \inst_midgetv_core.B_31\ : std_logic;
signal \inst_midgetv_core.sa42\ : std_logic;
signal \inst_midgetv_core.inst_progressctrl.badalignment\ : std_logic;
signal \inst_midgetv_core.buserror\ : std_logic;
signal \CONSTANT_ZERO_NET\ : std_logic;
signal \inst_midgetv_core.sa15\ : std_logic;
signal \inst_midgetv_core.sa32\ : std_logic;
signal \inst_midgetv_core.inst_ucodepc.maybranch_N_253\ : std_logic;
signal \inst_midgetv_core.sa30\ : std_logic;
signal \inst_midgetv_core.sa37\ : std_logic;
signal \inst_midgetv_core.sa25\ : std_logic;
signal \ADR_O_3\ : std_logic;
signal \inst_midgetv_core.inst_wai.genblk1_preWai1\ : std_logic;
signal \inst_midgetv_core.s_alu_carryin_0\ : std_logic;
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_28\ : std_logic;
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_31\ : std_logic;
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_30\ : std_logic;
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_29\ : std_logic;
signal \inst_midgetv_core.s_alu_carryin_1\ : std_logic;
signal \inst_midgetv_core.sa24\ : std_logic;
signal \inst_midgetv_core.inst_progressctrl.blka_usedefault\ : std_logic;
signal \inst_midgetv_core.inst_progressctrl.blka_en\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.genblk1_d_0\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_1\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_0\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_2\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_1\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_3\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_2\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_4\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_3\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_4\ : std_logic;
signal \inst_midgetv_core.lastshift\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.genblk1_d_2\ : std_logic;
signal \inst_midgetv_core.B_1\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.genblk1_d_3\ : std_logic;
signal \inst_midgetv_core.bmask_2\ : std_logic;
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.we\ : std_logic;
signal \inst_midgetv_core.bmask_3\ : std_logic;
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.we\ : std_logic;
signal \inst_midgetv_core.bmask_1\ : std_logic;
signal \inst_midgetv_core.iwe\ : std_logic;
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.we\ : std_logic;
signal \inst_midgetv_core.s_shift_1\ : std_logic;
signal \inst_midgetv_core.B_0\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_0\ : std_logic;
signal \CLK_c\ : std_logic;
signal \inst_midgetv_core.s_shift_0\ : std_logic;
signal \inst_midgetv_core.inst_shiftcounter.genblk1_d_1\ : std_logic;
signal \inst_midgetv_core.sa23\ : std_logic;
signal \ACK_I\ : std_logic;
signal \inst_midgetv_core.sa34\ : std_logic;
signal \inst_midgetv_core.sa40\ : std_logic;
signal \inst_midgetv_core.sram_stb\ : std_logic;
signal \STB_O\ : std_logic;
signal \inst_midgetv_core.sa20\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_sel0h\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_sel0hack\ : std_logic;
signal \inst_midgetv_core.sa26\ : std_logic;
signal \inst_midgetv_core.sa27\ : std_logic;
signal \inst_midgetv_core.ADR_O_8\ : std_logic;
signal \inst_midgetv_core.Wai_6\ : std_logic;
signal \inst_midgetv_core.INSTR_21\ : std_logic;
signal \inst_midgetv_core.INSTR_16\ : std_logic;
signal \inst_midgetv_core.INSTR_18\ : std_logic;
signal \inst_midgetv_core.INSTR_23\ : std_logic;
signal \inst_midgetv_core.INSTR_24\ : std_logic;
signal \inst_midgetv_core.INSTR_19\ : std_logic;
signal \inst_midgetv_core.INSTR_20\ : std_logic;
signal \inst_midgetv_core.INSTR_15\ : std_logic;
signal \inst_midgetv_core.B_6\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_b4a\ : std_logic;
signal \inst_midgetv_core.Rai_4\ : std_logic;
signal \inst_midgetv_core.B_2\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_sel_0\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_b0a\ : std_logic;
signal \inst_midgetv_core.Rai_0\ : std_logic;
signal \inst_midgetv_core.B_3\ : std_logic;
signal \inst_midgetv_core.sa21\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_b1a\ : std_logic;
signal \inst_midgetv_core.Rai_1\ : std_logic;
signal \inst_midgetv_core.B_7\ : std_logic;
signal \inst_midgetv_core.Rai_5\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_sel_3\ : std_logic;
signal \inst_midgetv_core.B_5\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_b3a\ : std_logic;
signal \inst_midgetv_core.Rai_3\ : std_logic;
signal \inst_midgetv_core.INSTR_22\ : std_logic;
signal \inst_midgetv_core.INSTR_17\ : std_logic;
signal \inst_midgetv_core.B_4\ : std_logic;
signal \inst_midgetv_core.sa22\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_b2a\ : std_logic;
signal \inst_midgetv_core.Rai_2\ : std_logic;
signal \inst_midgetv_core.B_10\ : std_logic;
signal \inst_midgetv_core.Rai_8\ : std_logic;
signal \inst_midgetv_core.B_11\ : std_logic;
signal \inst_midgetv_core.Rai_9\ : std_logic;
signal \inst_midgetv_core.B_8\ : std_logic;
signal \inst_midgetv_core.Rai_6\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_ss1\ : std_logic;
signal \inst_midgetv_core.B_9\ : std_logic;
signal \inst_midgetv_core.inst_rai.genblk1_ss0\ : std_logic;
signal \inst_midgetv_core.Rai_7\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \LED1_wire\ : std_logic;
signal \LED2_wire\ : std_logic;
signal \LED3_wire\ : std_logic;
signal \LED4_wire\ : std_logic;
signal \RX_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \CLK_wire\ <= CLK;
    LED1 <= \LED1_wire\;
    LED2 <= \LED2_wire\;
    LED3 <= \LED3_wire\;
    LED4 <= \LED4_wire\;
    \RX_wire\ <= RX;
    TX <= \TX_wire\;
    \DAT_O_3\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(13);
    \DAT_O_2\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(9);
    \DAT_O_1\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(5);
    \DAT_O_0\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(1);
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\ <= '0'&\N__13978\&\N__14113\&\N__14851\&\N__14947\&\N__14527\&\N__14755\&\N__13894\&\N__14251\&\N__15256\&\N__15043\;
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\ <= '0'&\N__10519\&\N__9667\&\N__11707\&\N__4696\&\N__6388\&\N__13237\&\N__10108\&\N__10210\&\N__10333\&\N__10426\;
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\ <= '0'&'0'&\N__14061\&'0'&'0'&'0'&\N__14195\&'0'&'0'&'0'&\N__12738\&'0'&'0'&'0'&\N__12493\&'0';
    \inst_midgetv_core.DAT_O_7\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(13);
    \inst_midgetv_core.DAT_O_6\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(9);
    \inst_midgetv_core.DAT_O_5\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(5);
    \inst_midgetv_core.DAT_O_4\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(1);
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\ <= '0'&\N__13972\&\N__14107\&\N__14845\&\N__14941\&\N__14521\&\N__14749\&\N__13888\&\N__14245\&\N__15250\&\N__15037\;
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\ <= '0'&\N__10513\&\N__9661\&\N__11701\&\N__4690\&\N__6382\&\N__13231\&\N__10102\&\N__10204\&\N__10327\&\N__10420\;
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\ <= '0'&'0'&\N__13927\&'0'&'0'&'0'&\N__14301\&'0'&'0'&'0'&\N__15293\&'0'&'0'&'0'&\N__15133\&'0';
    \inst_midgetv_core.DAT_O_11\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(13);
    \inst_midgetv_core.DAT_O_10\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(9);
    \inst_midgetv_core.DAT_O_9\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(5);
    \inst_midgetv_core.DAT_O_8\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(1);
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\ <= '0'&\N__13966\&\N__14101\&\N__14839\&\N__14935\&\N__14515\&\N__14743\&\N__13882\&\N__14239\&\N__15244\&\N__15031\;
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\ <= '0'&\N__10507\&\N__9655\&\N__11695\&\N__4684\&\N__6376\&\N__13225\&\N__10096\&\N__10198\&\N__10321\&\N__10414\;
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\ <= '0'&'0'&\N__14893\&'0'&'0'&'0'&\N__14988\&'0'&'0'&'0'&\N__14623\&'0'&'0'&'0'&\N__14796\&'0';
    \inst_midgetv_core.DAT_O_15\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(13);
    \inst_midgetv_core.DAT_O_14\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(9);
    \inst_midgetv_core.DAT_O_13\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(5);
    \inst_midgetv_core.DAT_O_12\ <= \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(1);
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\ <= '0'&\N__13960\&\N__14095\&\N__14833\&\N__14929\&\N__14509\&\N__14737\&\N__13876\&\N__14233\&\N__15238\&\N__15025\;
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\ <= '0'&\N__10501\&\N__9649\&\N__11689\&\N__4678\&\N__6370\&\N__13219\&\N__10090\&\N__10192\&\N__10315\&\N__10408\;
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\ <= '0'&'0'&\N__5587\&'0'&'0'&'0'&\N__5614\&'0'&'0'&'0'&\N__5641\&'0'&'0'&'0'&\N__5317\&'0';
    \inst_midgetv_core.DAT_O_19\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(13);
    \inst_midgetv_core.DAT_O_18\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(9);
    \inst_midgetv_core.DAT_O_17\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(5);
    \inst_midgetv_core.DAT_O_16\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(1);
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\ <= '0'&\N__13954\&\N__14089\&\N__14827\&\N__14923\&\N__14503\&\N__14731\&\N__13870\&\N__14227\&\N__15232\&\N__15019\;
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\ <= '0'&\N__10495\&\N__9643\&\N__11683\&\N__4672\&\N__6364\&\N__13213\&\N__10084\&\N__10186\&\N__10309\&\N__10402\;
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\ <= '0'&'0'&\N__5392\&'0'&'0'&'0'&\N__5499\&'0'&'0'&'0'&\N__5533\&'0'&'0'&'0'&\N__5563\&'0';
    \inst_midgetv_core.DAT_O_23\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(13);
    \inst_midgetv_core.DAT_O_22\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(9);
    \inst_midgetv_core.DAT_O_21\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(5);
    \inst_midgetv_core.DAT_O_20\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(1);
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\ <= '0'&\N__13948\&\N__14083\&\N__14821\&\N__14917\&\N__14497\&\N__14725\&\N__13864\&\N__14221\&\N__15226\&\N__15013\;
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\ <= '0'&\N__10489\&\N__9637\&\N__11677\&\N__4666\&\N__6358\&\N__13207\&\N__10078\&\N__10180\&\N__10303\&\N__10396\;
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\ <= '0'&'0'&\N__5827\&'0'&'0'&'0'&\N__5854\&'0'&'0'&'0'&\N__5887\&'0'&'0'&'0'&\N__5362\&'0';
    \inst_midgetv_core.DAT_O_27\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(13);
    \inst_midgetv_core.DAT_O_26\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(9);
    \inst_midgetv_core.DAT_O_25\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(5);
    \inst_midgetv_core.DAT_O_24\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\(1);
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\ <= '0'&\N__13942\&\N__14077\&\N__14815\&\N__14911\&\N__14491\&\N__14719\&\N__13858\&\N__14215\&\N__15220\&\N__15007\;
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\ <= '0'&\N__10483\&\N__9631\&\N__11671\&\N__4660\&\N__6352\&\N__13201\&\N__10072\&\N__10174\&\N__10297\&\N__10390\;
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\ <= '0'&'0'&\N__5701\&'0'&'0'&'0'&\N__5731\&'0'&'0'&'0'&\N__5761\&'0'&'0'&'0'&\N__5797\&'0';
    \DAT_O_31\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(13);
    \inst_midgetv_core.DAT_O_30\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(9);
    \inst_midgetv_core.DAT_O_29\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(5);
    \inst_midgetv_core.DAT_O_28\ <= \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\(1);
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\ <= '0'&\N__13936\&\N__14071\&\N__14809\&\N__14905\&\N__14485\&\N__14713\&\N__13852\&\N__14209\&\N__15214\&\N__15001\;
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\ <= '0'&\N__10477\&\N__9625\&\N__11665\&\N__4654\&\N__6346\&\N__13195\&\N__10066\&\N__10168\&\N__10291\&\N__10384\;
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\ <= '0'&'0'&\N__11434\&'0'&'0'&'0'&\N__8950\&'0'&'0'&'0'&\N__6202\&'0'&'0'&'0'&\N__5671\&'0';
    \inst_midgetv_core.sa20\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(15);
    \inst_midgetv_core.s_shift_1\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(14);
    \inst_midgetv_core.s_cyclecnt_1\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(13);
    \inst_midgetv_core.sa15\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(12);
    \inst_midgetv_core.sa14\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(11);
    \inst_midgetv_core.s_alu_2\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(10);
    \inst_midgetv_core.s_alu_1\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(9);
    \inst_midgetv_core.s_alu_0\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(8);
    \inst_midgetv_core.rinx_7\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(7);
    \inst_midgetv_core.rinx_6\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(6);
    \inst_midgetv_core.rinx_5\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(5);
    \inst_midgetv_core.rinx_4\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(4);
    \inst_midgetv_core.rinx_3\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(3);
    \inst_midgetv_core.rinx_2\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(2);
    \inst_midgetv_core.rinx_1\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(1);
    \inst_midgetv_core.rinx_0\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\(0);
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__7951\&\N__7795\&\N__7996\&\N__6268\&\N__7909\&\N__6226\&\N__8038\&\N__6325\;
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_31\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(15);
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_30\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(14);
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_29\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(13);
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_28\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(12);
    \inst_midgetv_core.sa43\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(11);
    \inst_midgetv_core.sa42\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(10);
    \inst_midgetv_core.sa41\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(9);
    \inst_midgetv_core.sa27\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(6);
    \inst_midgetv_core.sa26\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(5);
    \inst_midgetv_core.sa25\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(4);
    \inst_midgetv_core.sa24\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(3);
    \inst_midgetv_core.sa23\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(2);
    \inst_midgetv_core.sa22\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(1);
    \inst_midgetv_core.sa21\ <= \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\(0);
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__7944\&\N__7789\&\N__7990\&\N__6262\&\N__7903\&\N__6220\&\N__8032\&\N__6319\;
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';

    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100011101110000000011111111000000001111111110001000111111110000000011111111000000001111111100000000111111110110010011101110",
            INIT_0 => "1100110011001100000000000000000010001000111111110000100011001100000000000000000010111001100110011111111011101110010000000000000000001000111111110000000011111111000000001111111100000000111111110000000011111111000000011000100000000000100010000110010001000000"
        )
    port map (
            RDATA => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\,
            RADDR => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\,
            WADDR => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\,
            MASK => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_MASK_wire\,
            WDATA => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13823\,
            RE => \N__13008\,
            WCLKE => \N__9942\,
            WCLK => \N__13824\,
            WE => \N__13012\
        );

    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100011100011000000000011111011000101010000000111001110101000001010101010010001100010101010001000100010100000000010011000000",
            INIT_0 => "1100110011001100000000000000000001101100110100101100000010001100000000000000000010111011100110011101111111101110000000000000000001011100110000111111110111110000010001000100000101110000110011110100010011000001100000000000110000000000000000010100000001000100"
        )
    port map (
            RDATA => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\,
            RADDR => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\,
            WADDR => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\,
            MASK => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_MASK_wire\,
            WDATA => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13820\,
            RE => \N__13011\,
            WCLKE => \N__9943\,
            WCLK => \N__13821\,
            WE => \N__12978\
        );

    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000011110000111001000101111000100010101001101000101011110011000000101011011110001000100111110100000100000000000",
            INIT_0 => "1100110011001100000000000000000001000100010100000000000000000110000000000000000010011001100110011010101010101010000000000000010001000100011000000010011101100010010011100101000100000000111011100100111011010000000000000000000000000000000000000100000001000000"
        )
    port map (
            RDATA => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\,
            RADDR => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\,
            WADDR => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\,
            MASK => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_MASK_wire\,
            WDATA => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13816\,
            RE => \N__12905\,
            WCLKE => \N__12561\,
            WCLK => \N__13817\,
            WE => \N__12965\
        );

    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100011001000000001000001010100100000101000010001000101010001000000010000001100000001010000010110000101101001100010011000100",
            INIT_0 => "1100110011001100000000000000000010111100100110000100000000000000000000000000000010001001100110011010101010101010000000000000000010100000000001000111000100010100100001011110000101011010100000100010000010100100000000000000000000000000000000000100000001000100"
        )
    port map (
            RDATA => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\,
            RADDR => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\,
            WADDR => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\,
            MASK => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_MASK_wire\,
            WDATA => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13804\,
            RE => \N__12863\,
            WCLKE => \N__12565\,
            WCLK => \N__13805\,
            WE => \N__12907\
        );

    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010101000000111100001111000010010010001010001100100111010000111000010001000011000001010100001011010001000100110001000100",
            INIT_0 => "1100110011001100000000000000000010001000100010000000000000000100000000000000000010011001100110010010001000100010000000000000000000000000000011110000000010010001000011000001000100000010110011100000011000000000000000000000000000000000000000000100010000000100"
        )
    port map (
            RDATA => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\,
            RADDR => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\,
            WADDR => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\,
            MASK => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_MASK_wire\,
            WDATA => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13795\,
            RE => \N__12927\,
            WCLKE => \N__12645\,
            WCLK => \N__13796\,
            WE => \N__12926\
        );

    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110100001101000100001111001011010101000000000010100110000011001010001000100010101001100000010010100001000100010000101010101100",
            INIT_0 => "1100110011001100000000000000000010101010001111110010000000000100000000000000000010011001100110010010001000100010000000000000000000000000000000000000011110101001101001100100010111000000010000110010000000000000100000000000000000000000000000000100000001000000"
        )
    port map (
            RDATA => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\,
            RADDR => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\,
            WADDR => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\,
            MASK => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_MASK_wire\,
            WDATA => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13787\,
            RE => \N__12928\,
            WCLKE => \N__12649\,
            WCLK => \N__13788\,
            WE => \N__12982\
        );

    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100010011001000100010001000100011000100010000010111001000100000011001100110010001100010001000001000100010000000110010000100010",
            INIT_0 => "1100110011001100000000000000000011101110111000100000000000000000000000000000000010011001100110010010001000100010000000000000000001000000010000001111111100110000011001000100000000000000000000001100010001000001000000000000000000000000000000000100010001000000"
        )
    port map (
            RDATA => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RDATA_wire\,
            RADDR => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_RADDR_wire\,
            WADDR => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WADDR_wire\,
            MASK => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_MASK_wire\,
            WDATA => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrb.genblk1_mem_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13783\,
            RE => \N__12984\,
            WCLKE => \N__12618\,
            WCLK => \N__13784\,
            WE => \N__12983\
        );

    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "1100110011001100000000000000000011001110111011100000101010000000000000000000000010011001100110010010001000100010000000000000000001000100010001001111111111111111010001000100010000000000000000000100010001000100000000100010000010000000000000000100010000000100",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000100010001000100001000100010001010011001100110010011001100110011000101010001000101000100010001000100010001000100"
        )
    port map (
            RDATA => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RDATA_wire\,
            RADDR => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_RADDR_wire\,
            WADDR => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WADDR_wire\,
            MASK => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_MASK_wire\,
            WDATA => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.genblk1_ebrh.genblk1_mem_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13780\,
            RE => \N__12985\,
            WCLKE => \N__12619\,
            WCLK => \N__13781\,
            WE => \N__13009\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_F => "0101000011000111010000000100011001010000011111100111011001001001011101100110101101111100010001010000000000000000011101100001001101110110101010110101110011111010011101101101101111111100000000000100100011011101010100001110011001110110000111100111100101110010",
            INIT_E => "1100110011011110010000001111111000000000000000001101000000010001111110100101011000000000000000000101110011000110000000000000000001110110000111101100110011011110010111001011000111111010000110100000000000000000000000000000000001111001000111010000000000000000",
            INIT_D => "1111011011110100111101101111010001110110111001010111011001001001011001001001001001010000100100010000000000000000011101100001001101110110101000010100000011111110000000000000000001100100100100100111011000011110011110010000011001110110110010010111110000110111",
            INIT_C => "0101000001001111010000001111111000000000000000001101000000100110011101101110011000000000000000000101110010100101000000000000000001110001110010111111101101000111011110100110111111110010111000010000000000000000000000000000000001110110111010010000000000000000",
            INIT_B => "1111100111000001111110010001111111101011110111100111011001001001111111011011010111111010000110100000000000000000011101100001001101011100101111010101110010011010011101101001111000000000000000000000000000000000110011001101111001000100100100100101110010110010",
            INIT_A => "0111110011000101010000000011111100000000000000000100000000111111011100011001101000000000000000001110010000110100000000000000000001111100011000011110111011010000011111001010111110100110001110100000000000000000000000000000000001011100101101101011110001011110",
            INIT_9 => "0110100111110010011110011001111100000000000000000000000000000000000000000000000011000100001101000100000011111110011101100001001101100110100100111111100110111011110111001001010011100101001101001111000110010101111000010011010001000100100100100111011000110100",
            INIT_8 => "0111110010101001010000001111111000000000000000001101000000101001011101001110011000000000000000000000000000000000000000000000000001100001011111110100010000110100111110011111000011111010001000010000000000000000000000000000000001100001011111011011110010000101",
            INIT_7 => "0110000101111101011100011001000011100001001101000111011001001001011011100011001001101001111100100000000000000000000000000000000001100100011111010111100001110111010000000111001111110001111101000111000101110110011110100001101001110110000111100111100110111010",
            INIT_6 => "0111110011001111000000000000000000000000000000000101000000110001011110010111101000000000000000000000000000000000000000000000000001100110100100110110100111110010010100001110111111111010001010110000000000000000000000000000000001110010111101110000000000000000",
            INIT_5 => "0110111011011010111110010111000011111101111110110111011001001001011011100011001011111001010111010000000000000000000000000000000001111000100010110111101101010111011101100001111001111001111010110110111011011010111110010101010001101110110110101111000111100110",
            INIT_4 => "0111110011100110010000001111111000000000000000000101000000110001011010011011000001111100011001100111110001001011011111000110011001110001100011110110000101000111011111000110010111111010001010110000000000000000000000000000000001111100000010111111110001010000",
            INIT_3 => "1010000100111010101000010011010101111001000000110111011001001001011011100011001001111001001111010000000000000000011101100001001101110001110101111111110100000011111110010011011011101001110111100110010010000001011101001000011011111000001010110111011011100110",
            INIT_2 => "0111011011100110000000000000000001110110111001100100000000111110011101000011000000111100100101100111100000100001001111001001011001111100000111010111000000100111010010000000010010100110001101010101000011100110000000000000000001110000111001101011110001010010",
            INIT_1 => "0111011010110111010111001101010001110111111001101110111010100110011011100011001001110011111001100111010001000001011101100001001111111100011101001100111011011110011110010001011001111100000101011111100000010100000000000000000001111000000110101111100010001011",
            INIT_0 => "0111011011100110010100000001000001110110111001100111100100000100011100111000011000111100010110101111100010001011001111000101101011111011000010010111101000000111010010000000010001110100111001100101000011100110111111001011111011111001110100101011110000000001"
        )
    port map (
            RDATA => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RDATA_wire\,
            RADDR => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_RADDR_wire\,
            WADDR => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_WADDR_wire\,
            MASK => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_MASK_wire\,
            WDATA => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13826\,
            RE => \N__9807\,
            WCLKE => \N__11919\,
            WCLK => \GNDG0\,
            WE => 'L'
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000100001000000100000011100000000001000010000001000000111001100000110000100000000010001110000001000000010000000000100011100000010000000100000001000000011000000100000000100000000001000010000001000000001001000101000011000010010000001010000011000000110",
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_F => "0000001000000001000000100000000100000010000000010000000001100011000000100000000001010010000001010100000000000000000000000110011100000000011110010101001000000000000000000111110100000000010111110000001000000000000000100000000100000000011111011100001000000101",
            INIT_E => "0111010001010110000000100000000001000000000000000000001000000111000000100000001101000000000000000000001000000110010000000000000000000000011111010111010001010110010100100000010100000010000001110100000000000000010000000000000000000010000000000100000000000000",
            INIT_D => "1110000001000101111100000100000100000000011111010000000001100011010100000111000100000010000001010100000000000000000000000110011100000000011111010000001000000000010000000000000001010001111100010000000001111101110000100000010100000000010000110101001000000001",
            INIT_C => "0110001000000011000000100000000001000000000000000000001000000111000000011111101001000000000000000000001000000011010000000000000000000000011010000000010001101110000000100000000000000000010001110100000000000000010000000000000000000000011001010100000000000000",
            INIT_B => "1001001000000101100100100000010110010100010101100000000001100011101000000110010100000010000000110100000000000000000000000110011100000010000001100101001000000101000000100000000001000000000000000100000000000000011101000101011000000001111100010101001000000101",
            INIT_A => "0101001000000000000000100000011101000000000000000000001000000111000000000110110101000000000000000101000111110100010000000000000000000010000000000011001000000101010100100000001101000010000001110100000000000000010000000000000001010010000001010010010001100110",
            INIT_9 => "0000000000001110000011100000111001000000000000000100000000000000010000000000000000000001111101000000001000000000000000000110011100000000011110010100000001100101010100100000010100000001111101000000000001101101000000000110110001010001111100010000000111111010",
            INIT_8 => "0101001000000101000000100000000001000000000000000000001000000111010100000010000101000000000000000100000000000000010000000000000000000000011011100101000000100110000100100000010100000010000001110100000000000000010000000000000000000000011011010000011000000110",
            INIT_7 => "0000000001111101000000000110100000000001111101000000000001100011001100100000000100000000000101100100000000000000010000000000000001010000011011010000001000000001000000100000000111100010000001010000000001111110000000100000001100000000011111011100001000000101",
            INIT_6 => "0101001000000000010000000000000001000000000000000000001000000111000011100001011001000000000000000100000000000000010000000000000000000000011110010000000000011111011000100000000100000010000001110100000000000000010000000000000001100000010000110100000000000000",
            INIT_5 => "0000000001111101000100100000010110100000011001010000000001100011001100100000000101000000011001010100000000000000010000000000000000000010000001000000001000000100000000000111110111000010000001010000000001111101000100100000010100000000011111011101000000100101",
            INIT_4 => "0101001000000101000000100000000001000000000000000000001000000111000000010001110100111110000001110101001000000000001111100000011100000000011111010000000001101101010100100000010100000010000001110100000000000000010000000000000001010010000000000011011000000110",
            INIT_3 => "0100001000000111010000100000011111000000001001010000000001100011001100100000000110110000001001010100000000000000000000000110011101100000011010001010000000100101010000000010010110010100010101100000000001111001000000000110000100000010000001111000000000100001",
            INIT_2 => "0000000000100001010000000000000000000000001000010000001000000111010100100000000000100000010001110000001000000111001000000100011100000010000000000000000001000111000000100000000101000010000001110000001000000001010000000000000000000000001000010010010001100110",
            INIT_1 => "0000000001100101010100100000010100000000001000010010001000000101001100100000000100000000001000010000000001000101000000000110011100110100010101100111010001010110011000100000011001010010000000010000001000000111010000000000000000000010000001110000001000000111"
        )
    port map (
            RDATA => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RDATA_wire\,
            RADDR => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_RADDR_wire\,
            WADDR => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_WADDR_wire\,
            MASK => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_MASK_wire\,
            WDATA => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.ucode1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13825\,
            RE => \N__9806\,
            WCLKE => \N__11926\,
            WCLK => \GNDG0\,
            WE => 'L'
        );

    \CLK_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__15398\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15400\,
            DIN => \N__15399\,
            DOUT => \N__15398\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__15400\,
            PADOUT => \N__15399\,
            PADIN => \N__15398\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15389\,
            DIN => \N__15388\,
            DOUT => \N__15387\,
            PACKAGEPIN => \LED1_wire\
        );

    \LED1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__15389\,
            PADOUT => \N__15388\,
            PADIN => \N__15387\,
            CLOCKENABLE => \N__11484\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__6634\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__13778\,
            OUTPUTENABLE => '0'
        );

    \LED2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15380\,
            DIN => \N__15379\,
            DOUT => \N__15378\,
            PACKAGEPIN => \LED2_wire\
        );

    \LED2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__15380\,
            PADOUT => \N__15379\,
            PADIN => \N__15378\,
            CLOCKENABLE => \N__11484\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__6550\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__13778\,
            OUTPUTENABLE => '0'
        );

    \LED3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15371\,
            DIN => \N__15370\,
            DOUT => \N__15369\,
            PACKAGEPIN => \LED3_wire\
        );

    \LED3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__15371\,
            PADOUT => \N__15370\,
            PADIN => \N__15369\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10540\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED4_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15362\,
            DIN => \N__15361\,
            DOUT => \N__15360\,
            PACKAGEPIN => \LED4_wire\
        );

    \LED4_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__15362\,
            PADOUT => \N__15361\,
            PADIN => \N__15360\,
            CLOCKENABLE => \N__11488\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__6861\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__13779\,
            OUTPUTENABLE => '0'
        );

    \RX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15353\,
            DIN => \N__15352\,
            DOUT => \N__15351\,
            PACKAGEPIN => \RX_wire\
        );

    \RX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__15353\,
            PADOUT => \N__15352\,
            PADIN => \N__15351\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \meta_usartRX\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => \N__13827\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15344\,
            DIN => \N__15343\,
            DOUT => \N__15342\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__15344\,
            PADOUT => \N__15343\,
            PADIN => \N__15342\,
            CLOCKENABLE => \N__11581\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__6633\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__13828\,
            OUTPUTENABLE => '0'
        );

    \I__3895\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15320\
        );

    \I__3894\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15315\
        );

    \I__3893\ : InMux
    port map (
            O => \N__15323\,
            I => \N__15315\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__15320\,
            I => \N__15310\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__15315\,
            I => \N__15310\
        );

    \I__3890\ : Odrv12
    port map (
            O => \N__15310\,
            I => \inst_midgetv_core.inst_rai.genblk1_sel_3\
        );

    \I__3889\ : InMux
    port map (
            O => \N__15307\,
            I => \N__15303\
        );

    \I__3888\ : InMux
    port map (
            O => \N__15306\,
            I => \N__15300\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__15303\,
            I => \N__15297\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__15300\,
            I => \N__15294\
        );

    \I__3885\ : Span4Mux_v
    port map (
            O => \N__15297\,
            I => \N__15290\
        );

    \I__3884\ : Span4Mux_h
    port map (
            O => \N__15294\,
            I => \N__15287\
        );

    \I__3883\ : InMux
    port map (
            O => \N__15293\,
            I => \N__15284\
        );

    \I__3882\ : Sp12to4
    port map (
            O => \N__15290\,
            I => \N__15281\
        );

    \I__3881\ : Span4Mux_v
    port map (
            O => \N__15287\,
            I => \N__15278\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__15284\,
            I => \N__15275\
        );

    \I__3879\ : Span12Mux_h
    port map (
            O => \N__15281\,
            I => \N__15272\
        );

    \I__3878\ : Span4Mux_h
    port map (
            O => \N__15278\,
            I => \N__15269\
        );

    \I__3877\ : Odrv12
    port map (
            O => \N__15275\,
            I => \inst_midgetv_core.B_5\
        );

    \I__3876\ : Odrv12
    port map (
            O => \N__15272\,
            I => \inst_midgetv_core.B_5\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__15269\,
            I => \inst_midgetv_core.B_5\
        );

    \I__3874\ : InMux
    port map (
            O => \N__15262\,
            I => \N__15259\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__15259\,
            I => \inst_midgetv_core.inst_rai.genblk1_b3a\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__15256\,
            I => \N__15253\
        );

    \I__3871\ : CascadeBuf
    port map (
            O => \N__15253\,
            I => \N__15250\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__15250\,
            I => \N__15247\
        );

    \I__3869\ : CascadeBuf
    port map (
            O => \N__15247\,
            I => \N__15244\
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__15244\,
            I => \N__15241\
        );

    \I__3867\ : CascadeBuf
    port map (
            O => \N__15241\,
            I => \N__15238\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__15238\,
            I => \N__15235\
        );

    \I__3865\ : CascadeBuf
    port map (
            O => \N__15235\,
            I => \N__15232\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__15232\,
            I => \N__15229\
        );

    \I__3863\ : CascadeBuf
    port map (
            O => \N__15229\,
            I => \N__15226\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__15226\,
            I => \N__15223\
        );

    \I__3861\ : CascadeBuf
    port map (
            O => \N__15223\,
            I => \N__15220\
        );

    \I__3860\ : CascadeMux
    port map (
            O => \N__15220\,
            I => \N__15217\
        );

    \I__3859\ : CascadeBuf
    port map (
            O => \N__15217\,
            I => \N__15214\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__15214\,
            I => \N__15211\
        );

    \I__3857\ : InMux
    port map (
            O => \N__15211\,
            I => \N__15208\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__15208\,
            I => \inst_midgetv_core.Rai_3\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__15205\,
            I => \N__15202\
        );

    \I__3854\ : InMux
    port map (
            O => \N__15202\,
            I => \N__15199\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__15199\,
            I => \N__15194\
        );

    \I__3852\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15191\
        );

    \I__3851\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15188\
        );

    \I__3850\ : Span4Mux_s2_v
    port map (
            O => \N__15194\,
            I => \N__15185\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__15191\,
            I => \N__15180\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__15188\,
            I => \N__15180\
        );

    \I__3847\ : Span4Mux_v
    port map (
            O => \N__15185\,
            I => \N__15177\
        );

    \I__3846\ : Span12Mux_v
    port map (
            O => \N__15180\,
            I => \N__15174\
        );

    \I__3845\ : Span4Mux_v
    port map (
            O => \N__15177\,
            I => \N__15171\
        );

    \I__3844\ : Odrv12
    port map (
            O => \N__15174\,
            I => \inst_midgetv_core.INSTR_22\
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__15171\,
            I => \inst_midgetv_core.INSTR_22\
        );

    \I__3842\ : InMux
    port map (
            O => \N__15166\,
            I => \N__15163\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__15163\,
            I => \N__15159\
        );

    \I__3840\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15156\
        );

    \I__3839\ : Span4Mux_h
    port map (
            O => \N__15159\,
            I => \N__15153\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__15156\,
            I => \N__15150\
        );

    \I__3837\ : Span4Mux_v
    port map (
            O => \N__15153\,
            I => \N__15147\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__15150\,
            I => \N__15141\
        );

    \I__3835\ : Span4Mux_v
    port map (
            O => \N__15147\,
            I => \N__15141\
        );

    \I__3834\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15138\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__15141\,
            I => \inst_midgetv_core.INSTR_17\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__15138\,
            I => \inst_midgetv_core.INSTR_17\
        );

    \I__3831\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15128\
        );

    \I__3830\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15124\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__15131\,
            I => \N__15121\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__15128\,
            I => \N__15118\
        );

    \I__3827\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15115\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__15124\,
            I => \N__15112\
        );

    \I__3825\ : InMux
    port map (
            O => \N__15121\,
            I => \N__15109\
        );

    \I__3824\ : Span4Mux_v
    port map (
            O => \N__15118\,
            I => \N__15106\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__15115\,
            I => \N__15103\
        );

    \I__3822\ : Span12Mux_h
    port map (
            O => \N__15112\,
            I => \N__15100\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__15109\,
            I => \N__15097\
        );

    \I__3820\ : Sp12to4
    port map (
            O => \N__15106\,
            I => \N__15090\
        );

    \I__3819\ : Sp12to4
    port map (
            O => \N__15103\,
            I => \N__15090\
        );

    \I__3818\ : Span12Mux_v
    port map (
            O => \N__15100\,
            I => \N__15090\
        );

    \I__3817\ : Span4Mux_v
    port map (
            O => \N__15097\,
            I => \N__15087\
        );

    \I__3816\ : Odrv12
    port map (
            O => \N__15090\,
            I => \inst_midgetv_core.B_4\
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__15087\,
            I => \inst_midgetv_core.B_4\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__15082\,
            I => \N__15079\
        );

    \I__3813\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15074\
        );

    \I__3812\ : InMux
    port map (
            O => \N__15078\,
            I => \N__15069\
        );

    \I__3811\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15069\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__15074\,
            I => \N__15066\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__15069\,
            I => \N__15063\
        );

    \I__3808\ : Span4Mux_v
    port map (
            O => \N__15066\,
            I => \N__15058\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__15063\,
            I => \N__15058\
        );

    \I__3806\ : Span4Mux_v
    port map (
            O => \N__15058\,
            I => \N__15055\
        );

    \I__3805\ : Span4Mux_v
    port map (
            O => \N__15055\,
            I => \N__15052\
        );

    \I__3804\ : Odrv4
    port map (
            O => \N__15052\,
            I => \inst_midgetv_core.sa22\
        );

    \I__3803\ : InMux
    port map (
            O => \N__15049\,
            I => \N__15046\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__15046\,
            I => \inst_midgetv_core.inst_rai.genblk1_b2a\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__15043\,
            I => \N__15040\
        );

    \I__3800\ : CascadeBuf
    port map (
            O => \N__15040\,
            I => \N__15037\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__15037\,
            I => \N__15034\
        );

    \I__3798\ : CascadeBuf
    port map (
            O => \N__15034\,
            I => \N__15031\
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__15031\,
            I => \N__15028\
        );

    \I__3796\ : CascadeBuf
    port map (
            O => \N__15028\,
            I => \N__15025\
        );

    \I__3795\ : CascadeMux
    port map (
            O => \N__15025\,
            I => \N__15022\
        );

    \I__3794\ : CascadeBuf
    port map (
            O => \N__15022\,
            I => \N__15019\
        );

    \I__3793\ : CascadeMux
    port map (
            O => \N__15019\,
            I => \N__15016\
        );

    \I__3792\ : CascadeBuf
    port map (
            O => \N__15016\,
            I => \N__15013\
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__15013\,
            I => \N__15010\
        );

    \I__3790\ : CascadeBuf
    port map (
            O => \N__15010\,
            I => \N__15007\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__15007\,
            I => \N__15004\
        );

    \I__3788\ : CascadeBuf
    port map (
            O => \N__15004\,
            I => \N__15001\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__15001\,
            I => \N__14998\
        );

    \I__3786\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14995\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__14995\,
            I => \inst_midgetv_core.Rai_2\
        );

    \I__3784\ : InMux
    port map (
            O => \N__14992\,
            I => \N__14989\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__14989\,
            I => \N__14985\
        );

    \I__3782\ : InMux
    port map (
            O => \N__14988\,
            I => \N__14982\
        );

    \I__3781\ : Span4Mux_s1_v
    port map (
            O => \N__14985\,
            I => \N__14979\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__14982\,
            I => \N__14975\
        );

    \I__3779\ : Span4Mux_h
    port map (
            O => \N__14979\,
            I => \N__14972\
        );

    \I__3778\ : InMux
    port map (
            O => \N__14978\,
            I => \N__14969\
        );

    \I__3777\ : Span4Mux_v
    port map (
            O => \N__14975\,
            I => \N__14966\
        );

    \I__3776\ : Span4Mux_v
    port map (
            O => \N__14972\,
            I => \N__14963\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__14969\,
            I => \N__14960\
        );

    \I__3774\ : Span4Mux_h
    port map (
            O => \N__14966\,
            I => \N__14957\
        );

    \I__3773\ : Span4Mux_v
    port map (
            O => \N__14963\,
            I => \N__14952\
        );

    \I__3772\ : Span4Mux_v
    port map (
            O => \N__14960\,
            I => \N__14952\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__14957\,
            I => \inst_midgetv_core.B_10\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__14952\,
            I => \inst_midgetv_core.B_10\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__14947\,
            I => \N__14944\
        );

    \I__3768\ : CascadeBuf
    port map (
            O => \N__14944\,
            I => \N__14941\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__14941\,
            I => \N__14938\
        );

    \I__3766\ : CascadeBuf
    port map (
            O => \N__14938\,
            I => \N__14935\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__14935\,
            I => \N__14932\
        );

    \I__3764\ : CascadeBuf
    port map (
            O => \N__14932\,
            I => \N__14929\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__14929\,
            I => \N__14926\
        );

    \I__3762\ : CascadeBuf
    port map (
            O => \N__14926\,
            I => \N__14923\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__14923\,
            I => \N__14920\
        );

    \I__3760\ : CascadeBuf
    port map (
            O => \N__14920\,
            I => \N__14917\
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__14917\,
            I => \N__14914\
        );

    \I__3758\ : CascadeBuf
    port map (
            O => \N__14914\,
            I => \N__14911\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__14911\,
            I => \N__14908\
        );

    \I__3756\ : CascadeBuf
    port map (
            O => \N__14908\,
            I => \N__14905\
        );

    \I__3755\ : CascadeMux
    port map (
            O => \N__14905\,
            I => \N__14902\
        );

    \I__3754\ : InMux
    port map (
            O => \N__14902\,
            I => \N__14899\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__14899\,
            I => \N__14896\
        );

    \I__3752\ : Odrv4
    port map (
            O => \N__14896\,
            I => \inst_midgetv_core.Rai_8\
        );

    \I__3751\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14889\
        );

    \I__3750\ : InMux
    port map (
            O => \N__14892\,
            I => \N__14886\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__14889\,
            I => \N__14882\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__14886\,
            I => \N__14879\
        );

    \I__3747\ : InMux
    port map (
            O => \N__14885\,
            I => \N__14876\
        );

    \I__3746\ : Span4Mux_v
    port map (
            O => \N__14882\,
            I => \N__14873\
        );

    \I__3745\ : Span12Mux_s10_h
    port map (
            O => \N__14879\,
            I => \N__14870\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__14876\,
            I => \N__14867\
        );

    \I__3743\ : Span4Mux_h
    port map (
            O => \N__14873\,
            I => \N__14864\
        );

    \I__3742\ : Span12Mux_v
    port map (
            O => \N__14870\,
            I => \N__14861\
        );

    \I__3741\ : Span4Mux_h
    port map (
            O => \N__14867\,
            I => \N__14858\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__14864\,
            I => \inst_midgetv_core.B_11\
        );

    \I__3739\ : Odrv12
    port map (
            O => \N__14861\,
            I => \inst_midgetv_core.B_11\
        );

    \I__3738\ : Odrv4
    port map (
            O => \N__14858\,
            I => \inst_midgetv_core.B_11\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__14851\,
            I => \N__14848\
        );

    \I__3736\ : CascadeBuf
    port map (
            O => \N__14848\,
            I => \N__14845\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__14845\,
            I => \N__14842\
        );

    \I__3734\ : CascadeBuf
    port map (
            O => \N__14842\,
            I => \N__14839\
        );

    \I__3733\ : CascadeMux
    port map (
            O => \N__14839\,
            I => \N__14836\
        );

    \I__3732\ : CascadeBuf
    port map (
            O => \N__14836\,
            I => \N__14833\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__14833\,
            I => \N__14830\
        );

    \I__3730\ : CascadeBuf
    port map (
            O => \N__14830\,
            I => \N__14827\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__14827\,
            I => \N__14824\
        );

    \I__3728\ : CascadeBuf
    port map (
            O => \N__14824\,
            I => \N__14821\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__14821\,
            I => \N__14818\
        );

    \I__3726\ : CascadeBuf
    port map (
            O => \N__14818\,
            I => \N__14815\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__14815\,
            I => \N__14812\
        );

    \I__3724\ : CascadeBuf
    port map (
            O => \N__14812\,
            I => \N__14809\
        );

    \I__3723\ : CascadeMux
    port map (
            O => \N__14809\,
            I => \N__14806\
        );

    \I__3722\ : InMux
    port map (
            O => \N__14806\,
            I => \N__14803\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__14803\,
            I => \N__14800\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__14800\,
            I => \inst_midgetv_core.Rai_9\
        );

    \I__3719\ : InMux
    port map (
            O => \N__14797\,
            I => \N__14793\
        );

    \I__3718\ : InMux
    port map (
            O => \N__14796\,
            I => \N__14790\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__14793\,
            I => \N__14787\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__14790\,
            I => \N__14784\
        );

    \I__3715\ : Span4Mux_h
    port map (
            O => \N__14787\,
            I => \N__14781\
        );

    \I__3714\ : Span4Mux_v
    port map (
            O => \N__14784\,
            I => \N__14777\
        );

    \I__3713\ : Span4Mux_h
    port map (
            O => \N__14781\,
            I => \N__14774\
        );

    \I__3712\ : InMux
    port map (
            O => \N__14780\,
            I => \N__14771\
        );

    \I__3711\ : Span4Mux_h
    port map (
            O => \N__14777\,
            I => \N__14768\
        );

    \I__3710\ : Sp12to4
    port map (
            O => \N__14774\,
            I => \N__14765\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__14771\,
            I => \N__14762\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__14768\,
            I => \inst_midgetv_core.B_8\
        );

    \I__3707\ : Odrv12
    port map (
            O => \N__14765\,
            I => \inst_midgetv_core.B_8\
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__14762\,
            I => \inst_midgetv_core.B_8\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__14755\,
            I => \N__14752\
        );

    \I__3704\ : CascadeBuf
    port map (
            O => \N__14752\,
            I => \N__14749\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__14749\,
            I => \N__14746\
        );

    \I__3702\ : CascadeBuf
    port map (
            O => \N__14746\,
            I => \N__14743\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__14743\,
            I => \N__14740\
        );

    \I__3700\ : CascadeBuf
    port map (
            O => \N__14740\,
            I => \N__14737\
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__14737\,
            I => \N__14734\
        );

    \I__3698\ : CascadeBuf
    port map (
            O => \N__14734\,
            I => \N__14731\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__14731\,
            I => \N__14728\
        );

    \I__3696\ : CascadeBuf
    port map (
            O => \N__14728\,
            I => \N__14725\
        );

    \I__3695\ : CascadeMux
    port map (
            O => \N__14725\,
            I => \N__14722\
        );

    \I__3694\ : CascadeBuf
    port map (
            O => \N__14722\,
            I => \N__14719\
        );

    \I__3693\ : CascadeMux
    port map (
            O => \N__14719\,
            I => \N__14716\
        );

    \I__3692\ : CascadeBuf
    port map (
            O => \N__14716\,
            I => \N__14713\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__14713\,
            I => \N__14710\
        );

    \I__3690\ : InMux
    port map (
            O => \N__14710\,
            I => \N__14707\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__14707\,
            I => \inst_midgetv_core.Rai_6\
        );

    \I__3688\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14698\
        );

    \I__3687\ : CascadeMux
    port map (
            O => \N__14703\,
            I => \N__14693\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__14702\,
            I => \N__14689\
        );

    \I__3685\ : InMux
    port map (
            O => \N__14701\,
            I => \N__14686\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__14698\,
            I => \N__14679\
        );

    \I__3683\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14668\
        );

    \I__3682\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14668\
        );

    \I__3681\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14668\
        );

    \I__3680\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14668\
        );

    \I__3679\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14668\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__14686\,
            I => \N__14665\
        );

    \I__3677\ : InMux
    port map (
            O => \N__14685\,
            I => \N__14660\
        );

    \I__3676\ : InMux
    port map (
            O => \N__14684\,
            I => \N__14660\
        );

    \I__3675\ : InMux
    port map (
            O => \N__14683\,
            I => \N__14655\
        );

    \I__3674\ : InMux
    port map (
            O => \N__14682\,
            I => \N__14655\
        );

    \I__3673\ : Span4Mux_h
    port map (
            O => \N__14679\,
            I => \N__14648\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__14668\,
            I => \N__14639\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__14665\,
            I => \N__14639\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__14660\,
            I => \N__14639\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__14655\,
            I => \N__14639\
        );

    \I__3668\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14630\
        );

    \I__3667\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14630\
        );

    \I__3666\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14630\
        );

    \I__3665\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14630\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__14648\,
            I => \inst_midgetv_core.inst_rai.genblk1_ss1\
        );

    \I__3663\ : Odrv4
    port map (
            O => \N__14639\,
            I => \inst_midgetv_core.inst_rai.genblk1_ss1\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__14630\,
            I => \inst_midgetv_core.inst_rai.genblk1_ss1\
        );

    \I__3661\ : InMux
    port map (
            O => \N__14623\,
            I => \N__14620\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__14620\,
            I => \N__14616\
        );

    \I__3659\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14613\
        );

    \I__3658\ : Span4Mux_h
    port map (
            O => \N__14616\,
            I => \N__14610\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__14613\,
            I => \N__14607\
        );

    \I__3656\ : Sp12to4
    port map (
            O => \N__14610\,
            I => \N__14601\
        );

    \I__3655\ : Span12Mux_s8_h
    port map (
            O => \N__14607\,
            I => \N__14601\
        );

    \I__3654\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14598\
        );

    \I__3653\ : Span12Mux_v
    port map (
            O => \N__14601\,
            I => \N__14595\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__14598\,
            I => \N__14592\
        );

    \I__3651\ : Odrv12
    port map (
            O => \N__14595\,
            I => \inst_midgetv_core.B_9\
        );

    \I__3650\ : Odrv4
    port map (
            O => \N__14592\,
            I => \inst_midgetv_core.B_9\
        );

    \I__3649\ : InMux
    port map (
            O => \N__14587\,
            I => \N__14583\
        );

    \I__3648\ : InMux
    port map (
            O => \N__14586\,
            I => \N__14580\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__14583\,
            I => \N__14573\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__14580\,
            I => \N__14566\
        );

    \I__3645\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14561\
        );

    \I__3644\ : InMux
    port map (
            O => \N__14578\,
            I => \N__14561\
        );

    \I__3643\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14558\
        );

    \I__3642\ : InMux
    port map (
            O => \N__14576\,
            I => \N__14555\
        );

    \I__3641\ : Span4Mux_h
    port map (
            O => \N__14573\,
            I => \N__14552\
        );

    \I__3640\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14543\
        );

    \I__3639\ : InMux
    port map (
            O => \N__14571\,
            I => \N__14543\
        );

    \I__3638\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14543\
        );

    \I__3637\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14543\
        );

    \I__3636\ : Span4Mux_h
    port map (
            O => \N__14566\,
            I => \N__14536\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__14561\,
            I => \N__14536\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__14558\,
            I => \N__14536\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__14555\,
            I => \inst_midgetv_core.inst_rai.genblk1_ss0\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__14552\,
            I => \inst_midgetv_core.inst_rai.genblk1_ss0\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__14543\,
            I => \inst_midgetv_core.inst_rai.genblk1_ss0\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__14536\,
            I => \inst_midgetv_core.inst_rai.genblk1_ss0\
        );

    \I__3629\ : CascadeMux
    port map (
            O => \N__14527\,
            I => \N__14524\
        );

    \I__3628\ : CascadeBuf
    port map (
            O => \N__14524\,
            I => \N__14521\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__14521\,
            I => \N__14518\
        );

    \I__3626\ : CascadeBuf
    port map (
            O => \N__14518\,
            I => \N__14515\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__14515\,
            I => \N__14512\
        );

    \I__3624\ : CascadeBuf
    port map (
            O => \N__14512\,
            I => \N__14509\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__14509\,
            I => \N__14506\
        );

    \I__3622\ : CascadeBuf
    port map (
            O => \N__14506\,
            I => \N__14503\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__14503\,
            I => \N__14500\
        );

    \I__3620\ : CascadeBuf
    port map (
            O => \N__14500\,
            I => \N__14497\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__14497\,
            I => \N__14494\
        );

    \I__3618\ : CascadeBuf
    port map (
            O => \N__14494\,
            I => \N__14491\
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__14491\,
            I => \N__14488\
        );

    \I__3616\ : CascadeBuf
    port map (
            O => \N__14488\,
            I => \N__14485\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__14485\,
            I => \N__14482\
        );

    \I__3614\ : InMux
    port map (
            O => \N__14482\,
            I => \N__14479\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__14479\,
            I => \inst_midgetv_core.Rai_7\
        );

    \I__3612\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14473\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__14473\,
            I => \N__14469\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__14472\,
            I => \N__14466\
        );

    \I__3609\ : Span4Mux_h
    port map (
            O => \N__14469\,
            I => \N__14462\
        );

    \I__3608\ : InMux
    port map (
            O => \N__14466\,
            I => \N__14459\
        );

    \I__3607\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14456\
        );

    \I__3606\ : Span4Mux_v
    port map (
            O => \N__14462\,
            I => \N__14453\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__14459\,
            I => \N__14450\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__14456\,
            I => \N__14447\
        );

    \I__3603\ : Span4Mux_v
    port map (
            O => \N__14453\,
            I => \N__14442\
        );

    \I__3602\ : Span4Mux_v
    port map (
            O => \N__14450\,
            I => \N__14442\
        );

    \I__3601\ : Span4Mux_h
    port map (
            O => \N__14447\,
            I => \N__14439\
        );

    \I__3600\ : Span4Mux_h
    port map (
            O => \N__14442\,
            I => \N__14436\
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__14439\,
            I => \inst_midgetv_core.INSTR_24\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__14436\,
            I => \inst_midgetv_core.INSTR_24\
        );

    \I__3597\ : InMux
    port map (
            O => \N__14431\,
            I => \N__14427\
        );

    \I__3596\ : InMux
    port map (
            O => \N__14430\,
            I => \N__14424\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__14427\,
            I => \N__14421\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__14424\,
            I => \N__14417\
        );

    \I__3593\ : Span4Mux_v
    port map (
            O => \N__14421\,
            I => \N__14414\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__14420\,
            I => \N__14411\
        );

    \I__3591\ : Span4Mux_h
    port map (
            O => \N__14417\,
            I => \N__14408\
        );

    \I__3590\ : Span4Mux_v
    port map (
            O => \N__14414\,
            I => \N__14405\
        );

    \I__3589\ : InMux
    port map (
            O => \N__14411\,
            I => \N__14402\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__14408\,
            I => \inst_midgetv_core.INSTR_19\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__14405\,
            I => \inst_midgetv_core.INSTR_19\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__14402\,
            I => \inst_midgetv_core.INSTR_19\
        );

    \I__3585\ : CascadeMux
    port map (
            O => \N__14395\,
            I => \N__14392\
        );

    \I__3584\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14387\
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__14391\,
            I => \N__14383\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__14390\,
            I => \N__14380\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__14387\,
            I => \N__14377\
        );

    \I__3580\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14374\
        );

    \I__3579\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14371\
        );

    \I__3578\ : InMux
    port map (
            O => \N__14380\,
            I => \N__14368\
        );

    \I__3577\ : Span4Mux_h
    port map (
            O => \N__14377\,
            I => \N__14365\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__14374\,
            I => \N__14362\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__14371\,
            I => \N__14359\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__14368\,
            I => \N__14356\
        );

    \I__3573\ : Span4Mux_v
    port map (
            O => \N__14365\,
            I => \N__14353\
        );

    \I__3572\ : Sp12to4
    port map (
            O => \N__14362\,
            I => \N__14350\
        );

    \I__3571\ : Span4Mux_h
    port map (
            O => \N__14359\,
            I => \N__14345\
        );

    \I__3570\ : Span4Mux_h
    port map (
            O => \N__14356\,
            I => \N__14345\
        );

    \I__3569\ : Span4Mux_v
    port map (
            O => \N__14353\,
            I => \N__14342\
        );

    \I__3568\ : Odrv12
    port map (
            O => \N__14350\,
            I => \inst_midgetv_core.INSTR_20\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__14345\,
            I => \inst_midgetv_core.INSTR_20\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__14342\,
            I => \inst_midgetv_core.INSTR_20\
        );

    \I__3565\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14331\
        );

    \I__3564\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14328\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__14331\,
            I => \N__14325\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__14328\,
            I => \N__14321\
        );

    \I__3561\ : Span4Mux_v
    port map (
            O => \N__14325\,
            I => \N__14318\
        );

    \I__3560\ : InMux
    port map (
            O => \N__14324\,
            I => \N__14315\
        );

    \I__3559\ : Span4Mux_v
    port map (
            O => \N__14321\,
            I => \N__14310\
        );

    \I__3558\ : Span4Mux_v
    port map (
            O => \N__14318\,
            I => \N__14310\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__14315\,
            I => \N__14307\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__14310\,
            I => \inst_midgetv_core.INSTR_15\
        );

    \I__3555\ : Odrv12
    port map (
            O => \N__14307\,
            I => \inst_midgetv_core.INSTR_15\
        );

    \I__3554\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14298\
        );

    \I__3553\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14295\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__14298\,
            I => \N__14292\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__14295\,
            I => \N__14288\
        );

    \I__3550\ : Span4Mux_h
    port map (
            O => \N__14292\,
            I => \N__14285\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__14291\,
            I => \N__14282\
        );

    \I__3548\ : Span4Mux_v
    port map (
            O => \N__14288\,
            I => \N__14279\
        );

    \I__3547\ : Span4Mux_h
    port map (
            O => \N__14285\,
            I => \N__14276\
        );

    \I__3546\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14273\
        );

    \I__3545\ : Span4Mux_h
    port map (
            O => \N__14279\,
            I => \N__14270\
        );

    \I__3544\ : Sp12to4
    port map (
            O => \N__14276\,
            I => \N__14267\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__14273\,
            I => \N__14264\
        );

    \I__3542\ : Odrv4
    port map (
            O => \N__14270\,
            I => \inst_midgetv_core.B_6\
        );

    \I__3541\ : Odrv12
    port map (
            O => \N__14267\,
            I => \inst_midgetv_core.B_6\
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__14264\,
            I => \inst_midgetv_core.B_6\
        );

    \I__3539\ : InMux
    port map (
            O => \N__14257\,
            I => \N__14254\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__14254\,
            I => \inst_midgetv_core.inst_rai.genblk1_b4a\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__14251\,
            I => \N__14248\
        );

    \I__3536\ : CascadeBuf
    port map (
            O => \N__14248\,
            I => \N__14245\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__14245\,
            I => \N__14242\
        );

    \I__3534\ : CascadeBuf
    port map (
            O => \N__14242\,
            I => \N__14239\
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__14239\,
            I => \N__14236\
        );

    \I__3532\ : CascadeBuf
    port map (
            O => \N__14236\,
            I => \N__14233\
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__14233\,
            I => \N__14230\
        );

    \I__3530\ : CascadeBuf
    port map (
            O => \N__14230\,
            I => \N__14227\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__14227\,
            I => \N__14224\
        );

    \I__3528\ : CascadeBuf
    port map (
            O => \N__14224\,
            I => \N__14221\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__14221\,
            I => \N__14218\
        );

    \I__3526\ : CascadeBuf
    port map (
            O => \N__14218\,
            I => \N__14215\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__14215\,
            I => \N__14212\
        );

    \I__3524\ : CascadeBuf
    port map (
            O => \N__14212\,
            I => \N__14209\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__14209\,
            I => \N__14206\
        );

    \I__3522\ : InMux
    port map (
            O => \N__14206\,
            I => \N__14203\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__14203\,
            I => \inst_midgetv_core.Rai_4\
        );

    \I__3520\ : CascadeMux
    port map (
            O => \N__14200\,
            I => \N__14196\
        );

    \I__3519\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14191\
        );

    \I__3518\ : InMux
    port map (
            O => \N__14196\,
            I => \N__14188\
        );

    \I__3517\ : InMux
    port map (
            O => \N__14195\,
            I => \N__14185\
        );

    \I__3516\ : InMux
    port map (
            O => \N__14194\,
            I => \N__14182\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__14191\,
            I => \N__14179\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__14188\,
            I => \N__14176\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__14185\,
            I => \N__14173\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__14182\,
            I => \N__14170\
        );

    \I__3511\ : Span4Mux_v
    port map (
            O => \N__14179\,
            I => \N__14167\
        );

    \I__3510\ : Span4Mux_v
    port map (
            O => \N__14176\,
            I => \N__14164\
        );

    \I__3509\ : Span4Mux_v
    port map (
            O => \N__14173\,
            I => \N__14161\
        );

    \I__3508\ : Span4Mux_v
    port map (
            O => \N__14170\,
            I => \N__14158\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__14167\,
            I => \N__14155\
        );

    \I__3506\ : Span4Mux_h
    port map (
            O => \N__14164\,
            I => \N__14152\
        );

    \I__3505\ : Sp12to4
    port map (
            O => \N__14161\,
            I => \N__14149\
        );

    \I__3504\ : Span4Mux_h
    port map (
            O => \N__14158\,
            I => \N__14142\
        );

    \I__3503\ : Span4Mux_v
    port map (
            O => \N__14155\,
            I => \N__14142\
        );

    \I__3502\ : Span4Mux_v
    port map (
            O => \N__14152\,
            I => \N__14142\
        );

    \I__3501\ : Odrv12
    port map (
            O => \N__14149\,
            I => \inst_midgetv_core.B_2\
        );

    \I__3500\ : Odrv4
    port map (
            O => \N__14142\,
            I => \inst_midgetv_core.B_2\
        );

    \I__3499\ : InMux
    port map (
            O => \N__14137\,
            I => \N__14133\
        );

    \I__3498\ : InMux
    port map (
            O => \N__14136\,
            I => \N__14130\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__14133\,
            I => \N__14125\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__14130\,
            I => \N__14125\
        );

    \I__3495\ : Span12Mux_s5_v
    port map (
            O => \N__14125\,
            I => \N__14122\
        );

    \I__3494\ : Odrv12
    port map (
            O => \N__14122\,
            I => \inst_midgetv_core.inst_rai.genblk1_sel_0\
        );

    \I__3493\ : InMux
    port map (
            O => \N__14119\,
            I => \N__14116\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__14116\,
            I => \inst_midgetv_core.inst_rai.genblk1_b0a\
        );

    \I__3491\ : CascadeMux
    port map (
            O => \N__14113\,
            I => \N__14110\
        );

    \I__3490\ : CascadeBuf
    port map (
            O => \N__14110\,
            I => \N__14107\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__14107\,
            I => \N__14104\
        );

    \I__3488\ : CascadeBuf
    port map (
            O => \N__14104\,
            I => \N__14101\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__14101\,
            I => \N__14098\
        );

    \I__3486\ : CascadeBuf
    port map (
            O => \N__14098\,
            I => \N__14095\
        );

    \I__3485\ : CascadeMux
    port map (
            O => \N__14095\,
            I => \N__14092\
        );

    \I__3484\ : CascadeBuf
    port map (
            O => \N__14092\,
            I => \N__14089\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__14089\,
            I => \N__14086\
        );

    \I__3482\ : CascadeBuf
    port map (
            O => \N__14086\,
            I => \N__14083\
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__14083\,
            I => \N__14080\
        );

    \I__3480\ : CascadeBuf
    port map (
            O => \N__14080\,
            I => \N__14077\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__14077\,
            I => \N__14074\
        );

    \I__3478\ : CascadeBuf
    port map (
            O => \N__14074\,
            I => \N__14071\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__14071\,
            I => \N__14068\
        );

    \I__3476\ : InMux
    port map (
            O => \N__14068\,
            I => \N__14065\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__14065\,
            I => \inst_midgetv_core.Rai_0\
        );

    \I__3474\ : InMux
    port map (
            O => \N__14062\,
            I => \N__14058\
        );

    \I__3473\ : InMux
    port map (
            O => \N__14061\,
            I => \N__14055\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__14058\,
            I => \N__14052\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__14055\,
            I => \N__14048\
        );

    \I__3470\ : Span4Mux_v
    port map (
            O => \N__14052\,
            I => \N__14044\
        );

    \I__3469\ : InMux
    port map (
            O => \N__14051\,
            I => \N__14041\
        );

    \I__3468\ : Span4Mux_v
    port map (
            O => \N__14048\,
            I => \N__14038\
        );

    \I__3467\ : InMux
    port map (
            O => \N__14047\,
            I => \N__14035\
        );

    \I__3466\ : Span4Mux_h
    port map (
            O => \N__14044\,
            I => \N__14032\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__14041\,
            I => \N__14029\
        );

    \I__3464\ : Sp12to4
    port map (
            O => \N__14038\,
            I => \N__14024\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__14035\,
            I => \N__14024\
        );

    \I__3462\ : Span4Mux_v
    port map (
            O => \N__14032\,
            I => \N__14019\
        );

    \I__3461\ : Span4Mux_v
    port map (
            O => \N__14029\,
            I => \N__14019\
        );

    \I__3460\ : Odrv12
    port map (
            O => \N__14024\,
            I => \inst_midgetv_core.B_3\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__14019\,
            I => \inst_midgetv_core.B_3\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__14014\,
            I => \N__14011\
        );

    \I__3457\ : InMux
    port map (
            O => \N__14011\,
            I => \N__14008\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__14008\,
            I => \N__14004\
        );

    \I__3455\ : InMux
    port map (
            O => \N__14007\,
            I => \N__14001\
        );

    \I__3454\ : Span4Mux_h
    port map (
            O => \N__14004\,
            I => \N__13996\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__14001\,
            I => \N__13996\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__13996\,
            I => \N__13993\
        );

    \I__3451\ : Span4Mux_v
    port map (
            O => \N__13993\,
            I => \N__13990\
        );

    \I__3450\ : Span4Mux_v
    port map (
            O => \N__13990\,
            I => \N__13987\
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__13987\,
            I => \inst_midgetv_core.sa21\
        );

    \I__3448\ : InMux
    port map (
            O => \N__13984\,
            I => \N__13981\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__13981\,
            I => \inst_midgetv_core.inst_rai.genblk1_b1a\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__13978\,
            I => \N__13975\
        );

    \I__3445\ : CascadeBuf
    port map (
            O => \N__13975\,
            I => \N__13972\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__13972\,
            I => \N__13969\
        );

    \I__3443\ : CascadeBuf
    port map (
            O => \N__13969\,
            I => \N__13966\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__13966\,
            I => \N__13963\
        );

    \I__3441\ : CascadeBuf
    port map (
            O => \N__13963\,
            I => \N__13960\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__13960\,
            I => \N__13957\
        );

    \I__3439\ : CascadeBuf
    port map (
            O => \N__13957\,
            I => \N__13954\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__13954\,
            I => \N__13951\
        );

    \I__3437\ : CascadeBuf
    port map (
            O => \N__13951\,
            I => \N__13948\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__13948\,
            I => \N__13945\
        );

    \I__3435\ : CascadeBuf
    port map (
            O => \N__13945\,
            I => \N__13942\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__13942\,
            I => \N__13939\
        );

    \I__3433\ : CascadeBuf
    port map (
            O => \N__13939\,
            I => \N__13936\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__13936\,
            I => \N__13933\
        );

    \I__3431\ : InMux
    port map (
            O => \N__13933\,
            I => \N__13930\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__13930\,
            I => \inst_midgetv_core.Rai_1\
        );

    \I__3429\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13923\
        );

    \I__3428\ : InMux
    port map (
            O => \N__13926\,
            I => \N__13920\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__13923\,
            I => \N__13916\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__13920\,
            I => \N__13913\
        );

    \I__3425\ : InMux
    port map (
            O => \N__13919\,
            I => \N__13910\
        );

    \I__3424\ : Span12Mux_v
    port map (
            O => \N__13916\,
            I => \N__13907\
        );

    \I__3423\ : Span12Mux_h
    port map (
            O => \N__13913\,
            I => \N__13904\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__13910\,
            I => \N__13901\
        );

    \I__3421\ : Odrv12
    port map (
            O => \N__13907\,
            I => \inst_midgetv_core.B_7\
        );

    \I__3420\ : Odrv12
    port map (
            O => \N__13904\,
            I => \inst_midgetv_core.B_7\
        );

    \I__3419\ : Odrv4
    port map (
            O => \N__13901\,
            I => \inst_midgetv_core.B_7\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__13894\,
            I => \N__13891\
        );

    \I__3417\ : CascadeBuf
    port map (
            O => \N__13891\,
            I => \N__13888\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__13888\,
            I => \N__13885\
        );

    \I__3415\ : CascadeBuf
    port map (
            O => \N__13885\,
            I => \N__13882\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__13882\,
            I => \N__13879\
        );

    \I__3413\ : CascadeBuf
    port map (
            O => \N__13879\,
            I => \N__13876\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__13876\,
            I => \N__13873\
        );

    \I__3411\ : CascadeBuf
    port map (
            O => \N__13873\,
            I => \N__13870\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__13870\,
            I => \N__13867\
        );

    \I__3409\ : CascadeBuf
    port map (
            O => \N__13867\,
            I => \N__13864\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__13864\,
            I => \N__13861\
        );

    \I__3407\ : CascadeBuf
    port map (
            O => \N__13861\,
            I => \N__13858\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__13858\,
            I => \N__13855\
        );

    \I__3405\ : CascadeBuf
    port map (
            O => \N__13855\,
            I => \N__13852\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__13852\,
            I => \N__13849\
        );

    \I__3403\ : InMux
    port map (
            O => \N__13849\,
            I => \N__13846\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__13846\,
            I => \inst_midgetv_core.Rai_5\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__13843\,
            I => \N__13839\
        );

    \I__3400\ : InMux
    port map (
            O => \N__13842\,
            I => \N__13836\
        );

    \I__3399\ : InMux
    port map (
            O => \N__13839\,
            I => \N__13833\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__13836\,
            I => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_0\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__13833\,
            I => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_0\
        );

    \I__3396\ : ClkMux
    port map (
            O => \N__13828\,
            I => \N__13675\
        );

    \I__3395\ : ClkMux
    port map (
            O => \N__13827\,
            I => \N__13675\
        );

    \I__3394\ : ClkMux
    port map (
            O => \N__13826\,
            I => \N__13675\
        );

    \I__3393\ : ClkMux
    port map (
            O => \N__13825\,
            I => \N__13675\
        );

    \I__3392\ : ClkMux
    port map (
            O => \N__13824\,
            I => \N__13675\
        );

    \I__3391\ : ClkMux
    port map (
            O => \N__13823\,
            I => \N__13675\
        );

    \I__3390\ : ClkMux
    port map (
            O => \N__13822\,
            I => \N__13675\
        );

    \I__3389\ : ClkMux
    port map (
            O => \N__13821\,
            I => \N__13675\
        );

    \I__3388\ : ClkMux
    port map (
            O => \N__13820\,
            I => \N__13675\
        );

    \I__3387\ : ClkMux
    port map (
            O => \N__13819\,
            I => \N__13675\
        );

    \I__3386\ : ClkMux
    port map (
            O => \N__13818\,
            I => \N__13675\
        );

    \I__3385\ : ClkMux
    port map (
            O => \N__13817\,
            I => \N__13675\
        );

    \I__3384\ : ClkMux
    port map (
            O => \N__13816\,
            I => \N__13675\
        );

    \I__3383\ : ClkMux
    port map (
            O => \N__13815\,
            I => \N__13675\
        );

    \I__3382\ : ClkMux
    port map (
            O => \N__13814\,
            I => \N__13675\
        );

    \I__3381\ : ClkMux
    port map (
            O => \N__13813\,
            I => \N__13675\
        );

    \I__3380\ : ClkMux
    port map (
            O => \N__13812\,
            I => \N__13675\
        );

    \I__3379\ : ClkMux
    port map (
            O => \N__13811\,
            I => \N__13675\
        );

    \I__3378\ : ClkMux
    port map (
            O => \N__13810\,
            I => \N__13675\
        );

    \I__3377\ : ClkMux
    port map (
            O => \N__13809\,
            I => \N__13675\
        );

    \I__3376\ : ClkMux
    port map (
            O => \N__13808\,
            I => \N__13675\
        );

    \I__3375\ : ClkMux
    port map (
            O => \N__13807\,
            I => \N__13675\
        );

    \I__3374\ : ClkMux
    port map (
            O => \N__13806\,
            I => \N__13675\
        );

    \I__3373\ : ClkMux
    port map (
            O => \N__13805\,
            I => \N__13675\
        );

    \I__3372\ : ClkMux
    port map (
            O => \N__13804\,
            I => \N__13675\
        );

    \I__3371\ : ClkMux
    port map (
            O => \N__13803\,
            I => \N__13675\
        );

    \I__3370\ : ClkMux
    port map (
            O => \N__13802\,
            I => \N__13675\
        );

    \I__3369\ : ClkMux
    port map (
            O => \N__13801\,
            I => \N__13675\
        );

    \I__3368\ : ClkMux
    port map (
            O => \N__13800\,
            I => \N__13675\
        );

    \I__3367\ : ClkMux
    port map (
            O => \N__13799\,
            I => \N__13675\
        );

    \I__3366\ : ClkMux
    port map (
            O => \N__13798\,
            I => \N__13675\
        );

    \I__3365\ : ClkMux
    port map (
            O => \N__13797\,
            I => \N__13675\
        );

    \I__3364\ : ClkMux
    port map (
            O => \N__13796\,
            I => \N__13675\
        );

    \I__3363\ : ClkMux
    port map (
            O => \N__13795\,
            I => \N__13675\
        );

    \I__3362\ : ClkMux
    port map (
            O => \N__13794\,
            I => \N__13675\
        );

    \I__3361\ : ClkMux
    port map (
            O => \N__13793\,
            I => \N__13675\
        );

    \I__3360\ : ClkMux
    port map (
            O => \N__13792\,
            I => \N__13675\
        );

    \I__3359\ : ClkMux
    port map (
            O => \N__13791\,
            I => \N__13675\
        );

    \I__3358\ : ClkMux
    port map (
            O => \N__13790\,
            I => \N__13675\
        );

    \I__3357\ : ClkMux
    port map (
            O => \N__13789\,
            I => \N__13675\
        );

    \I__3356\ : ClkMux
    port map (
            O => \N__13788\,
            I => \N__13675\
        );

    \I__3355\ : ClkMux
    port map (
            O => \N__13787\,
            I => \N__13675\
        );

    \I__3354\ : ClkMux
    port map (
            O => \N__13786\,
            I => \N__13675\
        );

    \I__3353\ : ClkMux
    port map (
            O => \N__13785\,
            I => \N__13675\
        );

    \I__3352\ : ClkMux
    port map (
            O => \N__13784\,
            I => \N__13675\
        );

    \I__3351\ : ClkMux
    port map (
            O => \N__13783\,
            I => \N__13675\
        );

    \I__3350\ : ClkMux
    port map (
            O => \N__13782\,
            I => \N__13675\
        );

    \I__3349\ : ClkMux
    port map (
            O => \N__13781\,
            I => \N__13675\
        );

    \I__3348\ : ClkMux
    port map (
            O => \N__13780\,
            I => \N__13675\
        );

    \I__3347\ : ClkMux
    port map (
            O => \N__13779\,
            I => \N__13675\
        );

    \I__3346\ : ClkMux
    port map (
            O => \N__13778\,
            I => \N__13675\
        );

    \I__3345\ : GlobalMux
    port map (
            O => \N__13675\,
            I => \N__13672\
        );

    \I__3344\ : gio2CtrlBuf
    port map (
            O => \N__13672\,
            I => \CLK_c\
        );

    \I__3343\ : InMux
    port map (
            O => \N__13669\,
            I => \N__13661\
        );

    \I__3342\ : InMux
    port map (
            O => \N__13668\,
            I => \N__13661\
        );

    \I__3341\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13655\
        );

    \I__3340\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13655\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__13661\,
            I => \N__13652\
        );

    \I__3338\ : InMux
    port map (
            O => \N__13660\,
            I => \N__13649\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__13655\,
            I => \N__13646\
        );

    \I__3336\ : Span4Mux_h
    port map (
            O => \N__13652\,
            I => \N__13641\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__13649\,
            I => \N__13641\
        );

    \I__3334\ : Odrv12
    port map (
            O => \N__13646\,
            I => \inst_midgetv_core.s_shift_0\
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__13641\,
            I => \inst_midgetv_core.s_shift_0\
        );

    \I__3332\ : InMux
    port map (
            O => \N__13636\,
            I => \N__13633\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__13633\,
            I => \inst_midgetv_core.inst_shiftcounter.genblk1_d_1\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__13630\,
            I => \N__13627\
        );

    \I__3329\ : InMux
    port map (
            O => \N__13627\,
            I => \N__13624\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__13624\,
            I => \N__13621\
        );

    \I__3327\ : Span4Mux_v
    port map (
            O => \N__13621\,
            I => \N__13618\
        );

    \I__3326\ : Odrv4
    port map (
            O => \N__13618\,
            I => \inst_midgetv_core.sa23\
        );

    \I__3325\ : InMux
    port map (
            O => \N__13615\,
            I => \N__13612\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__13612\,
            I => \N__13609\
        );

    \I__3323\ : Span4Mux_h
    port map (
            O => \N__13609\,
            I => \N__13605\
        );

    \I__3322\ : InMux
    port map (
            O => \N__13608\,
            I => \N__13602\
        );

    \I__3321\ : Odrv4
    port map (
            O => \N__13605\,
            I => \ACK_I\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__13602\,
            I => \ACK_I\
        );

    \I__3319\ : InMux
    port map (
            O => \N__13597\,
            I => \N__13591\
        );

    \I__3318\ : InMux
    port map (
            O => \N__13596\,
            I => \N__13591\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__13591\,
            I => \N__13588\
        );

    \I__3316\ : Odrv12
    port map (
            O => \N__13588\,
            I => \inst_midgetv_core.sa34\
        );

    \I__3315\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13576\
        );

    \I__3314\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13576\
        );

    \I__3313\ : InMux
    port map (
            O => \N__13583\,
            I => \N__13576\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__13576\,
            I => \N__13573\
        );

    \I__3311\ : Odrv12
    port map (
            O => \N__13573\,
            I => \inst_midgetv_core.sa40\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__13570\,
            I => \N__13566\
        );

    \I__3309\ : InMux
    port map (
            O => \N__13569\,
            I => \N__13560\
        );

    \I__3308\ : InMux
    port map (
            O => \N__13566\,
            I => \N__13560\
        );

    \I__3307\ : InMux
    port map (
            O => \N__13565\,
            I => \N__13557\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__13560\,
            I => \N__13554\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__13557\,
            I => \inst_midgetv_core.sram_stb\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__13554\,
            I => \inst_midgetv_core.sram_stb\
        );

    \I__3303\ : InMux
    port map (
            O => \N__13549\,
            I => \N__13546\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__13546\,
            I => \N__13542\
        );

    \I__3301\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13539\
        );

    \I__3300\ : Span4Mux_v
    port map (
            O => \N__13542\,
            I => \N__13528\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__13539\,
            I => \N__13528\
        );

    \I__3298\ : InMux
    port map (
            O => \N__13538\,
            I => \N__13525\
        );

    \I__3297\ : InMux
    port map (
            O => \N__13537\,
            I => \N__13522\
        );

    \I__3296\ : InMux
    port map (
            O => \N__13536\,
            I => \N__13515\
        );

    \I__3295\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13515\
        );

    \I__3294\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13512\
        );

    \I__3293\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13509\
        );

    \I__3292\ : Span4Mux_h
    port map (
            O => \N__13528\,
            I => \N__13506\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__13525\,
            I => \N__13501\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__13522\,
            I => \N__13501\
        );

    \I__3289\ : InMux
    port map (
            O => \N__13521\,
            I => \N__13496\
        );

    \I__3288\ : InMux
    port map (
            O => \N__13520\,
            I => \N__13496\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__13515\,
            I => \N__13493\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__13512\,
            I => \N__13490\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__13509\,
            I => \STB_O\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__13506\,
            I => \STB_O\
        );

    \I__3283\ : Odrv12
    port map (
            O => \N__13501\,
            I => \STB_O\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__13496\,
            I => \STB_O\
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__13493\,
            I => \STB_O\
        );

    \I__3280\ : Odrv4
    port map (
            O => \N__13490\,
            I => \STB_O\
        );

    \I__3279\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13474\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__13474\,
            I => \N__13471\
        );

    \I__3277\ : Span4Mux_v
    port map (
            O => \N__13471\,
            I => \N__13468\
        );

    \I__3276\ : Span4Mux_v
    port map (
            O => \N__13468\,
            I => \N__13465\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__13465\,
            I => \inst_midgetv_core.sa20\
        );

    \I__3274\ : InMux
    port map (
            O => \N__13462\,
            I => \N__13459\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__13459\,
            I => \inst_midgetv_core.inst_rai.genblk1_sel0h\
        );

    \I__3272\ : InMux
    port map (
            O => \N__13456\,
            I => \N__13453\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__13453\,
            I => \inst_midgetv_core.inst_rai.genblk1_sel0hack\
        );

    \I__3270\ : InMux
    port map (
            O => \N__13450\,
            I => \N__13446\
        );

    \I__3269\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13443\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__13446\,
            I => \N__13436\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__13443\,
            I => \N__13436\
        );

    \I__3266\ : InMux
    port map (
            O => \N__13442\,
            I => \N__13433\
        );

    \I__3265\ : InMux
    port map (
            O => \N__13441\,
            I => \N__13427\
        );

    \I__3264\ : Span4Mux_h
    port map (
            O => \N__13436\,
            I => \N__13422\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__13433\,
            I => \N__13422\
        );

    \I__3262\ : CascadeMux
    port map (
            O => \N__13432\,
            I => \N__13418\
        );

    \I__3261\ : CascadeMux
    port map (
            O => \N__13431\,
            I => \N__13414\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__13430\,
            I => \N__13410\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__13427\,
            I => \N__13407\
        );

    \I__3258\ : Span4Mux_v
    port map (
            O => \N__13422\,
            I => \N__13404\
        );

    \I__3257\ : InMux
    port map (
            O => \N__13421\,
            I => \N__13391\
        );

    \I__3256\ : InMux
    port map (
            O => \N__13418\,
            I => \N__13391\
        );

    \I__3255\ : InMux
    port map (
            O => \N__13417\,
            I => \N__13391\
        );

    \I__3254\ : InMux
    port map (
            O => \N__13414\,
            I => \N__13391\
        );

    \I__3253\ : InMux
    port map (
            O => \N__13413\,
            I => \N__13391\
        );

    \I__3252\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13391\
        );

    \I__3251\ : Span4Mux_h
    port map (
            O => \N__13407\,
            I => \N__13387\
        );

    \I__3250\ : Span4Mux_v
    port map (
            O => \N__13404\,
            I => \N__13382\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__13391\,
            I => \N__13382\
        );

    \I__3248\ : InMux
    port map (
            O => \N__13390\,
            I => \N__13379\
        );

    \I__3247\ : Span4Mux_h
    port map (
            O => \N__13387\,
            I => \N__13376\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__13382\,
            I => \N__13373\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__13379\,
            I => \inst_midgetv_core.sa26\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__13376\,
            I => \inst_midgetv_core.sa26\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__13373\,
            I => \inst_midgetv_core.sa26\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__13366\,
            I => \N__13362\
        );

    \I__3241\ : CascadeMux
    port map (
            O => \N__13365\,
            I => \N__13358\
        );

    \I__3240\ : InMux
    port map (
            O => \N__13362\,
            I => \N__13354\
        );

    \I__3239\ : InMux
    port map (
            O => \N__13361\,
            I => \N__13351\
        );

    \I__3238\ : InMux
    port map (
            O => \N__13358\,
            I => \N__13348\
        );

    \I__3237\ : InMux
    port map (
            O => \N__13357\,
            I => \N__13345\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__13354\,
            I => \N__13339\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__13351\,
            I => \N__13339\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__13348\,
            I => \N__13336\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__13345\,
            I => \N__13333\
        );

    \I__3232\ : InMux
    port map (
            O => \N__13344\,
            I => \N__13324\
        );

    \I__3231\ : Span4Mux_h
    port map (
            O => \N__13339\,
            I => \N__13321\
        );

    \I__3230\ : Span4Mux_h
    port map (
            O => \N__13336\,
            I => \N__13316\
        );

    \I__3229\ : Span4Mux_v
    port map (
            O => \N__13333\,
            I => \N__13316\
        );

    \I__3228\ : InMux
    port map (
            O => \N__13332\,
            I => \N__13303\
        );

    \I__3227\ : InMux
    port map (
            O => \N__13331\,
            I => \N__13303\
        );

    \I__3226\ : InMux
    port map (
            O => \N__13330\,
            I => \N__13303\
        );

    \I__3225\ : InMux
    port map (
            O => \N__13329\,
            I => \N__13303\
        );

    \I__3224\ : InMux
    port map (
            O => \N__13328\,
            I => \N__13303\
        );

    \I__3223\ : InMux
    port map (
            O => \N__13327\,
            I => \N__13303\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__13324\,
            I => \N__13300\
        );

    \I__3221\ : Span4Mux_v
    port map (
            O => \N__13321\,
            I => \N__13291\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__13316\,
            I => \N__13291\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__13303\,
            I => \N__13291\
        );

    \I__3218\ : Span12Mux_v
    port map (
            O => \N__13300\,
            I => \N__13288\
        );

    \I__3217\ : InMux
    port map (
            O => \N__13299\,
            I => \N__13283\
        );

    \I__3216\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13283\
        );

    \I__3215\ : Span4Mux_h
    port map (
            O => \N__13291\,
            I => \N__13280\
        );

    \I__3214\ : Odrv12
    port map (
            O => \N__13288\,
            I => \inst_midgetv_core.sa27\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__13283\,
            I => \inst_midgetv_core.sa27\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__13280\,
            I => \inst_midgetv_core.sa27\
        );

    \I__3211\ : InMux
    port map (
            O => \N__13273\,
            I => \N__13270\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__13270\,
            I => \N__13267\
        );

    \I__3209\ : Span4Mux_v
    port map (
            O => \N__13267\,
            I => \N__13262\
        );

    \I__3208\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13259\
        );

    \I__3207\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13255\
        );

    \I__3206\ : Span4Mux_h
    port map (
            O => \N__13262\,
            I => \N__13250\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__13259\,
            I => \N__13250\
        );

    \I__3204\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13247\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__13255\,
            I => \N__13244\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__13250\,
            I => \inst_midgetv_core.ADR_O_8\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__13247\,
            I => \inst_midgetv_core.ADR_O_8\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__13244\,
            I => \inst_midgetv_core.ADR_O_8\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__13237\,
            I => \N__13234\
        );

    \I__3198\ : CascadeBuf
    port map (
            O => \N__13234\,
            I => \N__13231\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__13231\,
            I => \N__13228\
        );

    \I__3196\ : CascadeBuf
    port map (
            O => \N__13228\,
            I => \N__13225\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__13225\,
            I => \N__13222\
        );

    \I__3194\ : CascadeBuf
    port map (
            O => \N__13222\,
            I => \N__13219\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__13219\,
            I => \N__13216\
        );

    \I__3192\ : CascadeBuf
    port map (
            O => \N__13216\,
            I => \N__13213\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__13213\,
            I => \N__13210\
        );

    \I__3190\ : CascadeBuf
    port map (
            O => \N__13210\,
            I => \N__13207\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__13207\,
            I => \N__13204\
        );

    \I__3188\ : CascadeBuf
    port map (
            O => \N__13204\,
            I => \N__13201\
        );

    \I__3187\ : CascadeMux
    port map (
            O => \N__13201\,
            I => \N__13198\
        );

    \I__3186\ : CascadeBuf
    port map (
            O => \N__13198\,
            I => \N__13195\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__13195\,
            I => \N__13192\
        );

    \I__3184\ : InMux
    port map (
            O => \N__13192\,
            I => \N__13189\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__13189\,
            I => \N__13186\
        );

    \I__3182\ : Span12Mux_s11_v
    port map (
            O => \N__13186\,
            I => \N__13183\
        );

    \I__3181\ : Odrv12
    port map (
            O => \N__13183\,
            I => \inst_midgetv_core.Wai_6\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__13180\,
            I => \N__13177\
        );

    \I__3179\ : InMux
    port map (
            O => \N__13177\,
            I => \N__13173\
        );

    \I__3178\ : InMux
    port map (
            O => \N__13176\,
            I => \N__13170\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__13173\,
            I => \N__13166\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__13170\,
            I => \N__13163\
        );

    \I__3175\ : InMux
    port map (
            O => \N__13169\,
            I => \N__13160\
        );

    \I__3174\ : Span4Mux_v
    port map (
            O => \N__13166\,
            I => \N__13157\
        );

    \I__3173\ : Span4Mux_v
    port map (
            O => \N__13163\,
            I => \N__13154\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__13160\,
            I => \N__13151\
        );

    \I__3171\ : Span4Mux_v
    port map (
            O => \N__13157\,
            I => \N__13148\
        );

    \I__3170\ : Odrv4
    port map (
            O => \N__13154\,
            I => \inst_midgetv_core.INSTR_21\
        );

    \I__3169\ : Odrv12
    port map (
            O => \N__13151\,
            I => \inst_midgetv_core.INSTR_21\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__13148\,
            I => \inst_midgetv_core.INSTR_21\
        );

    \I__3167\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13138\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__13138\,
            I => \N__13134\
        );

    \I__3165\ : InMux
    port map (
            O => \N__13137\,
            I => \N__13131\
        );

    \I__3164\ : Span4Mux_h
    port map (
            O => \N__13134\,
            I => \N__13127\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__13131\,
            I => \N__13124\
        );

    \I__3162\ : InMux
    port map (
            O => \N__13130\,
            I => \N__13121\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__13127\,
            I => \N__13118\
        );

    \I__3160\ : Span12Mux_s11_v
    port map (
            O => \N__13124\,
            I => \N__13115\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__13121\,
            I => \N__13112\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__13118\,
            I => \inst_midgetv_core.INSTR_16\
        );

    \I__3157\ : Odrv12
    port map (
            O => \N__13115\,
            I => \inst_midgetv_core.INSTR_16\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__13112\,
            I => \inst_midgetv_core.INSTR_16\
        );

    \I__3155\ : CascadeMux
    port map (
            O => \N__13105\,
            I => \N__13101\
        );

    \I__3154\ : InMux
    port map (
            O => \N__13104\,
            I => \N__13098\
        );

    \I__3153\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13095\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__13098\,
            I => \N__13091\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__13095\,
            I => \N__13088\
        );

    \I__3150\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13085\
        );

    \I__3149\ : Span4Mux_v
    port map (
            O => \N__13091\,
            I => \N__13082\
        );

    \I__3148\ : Span4Mux_v
    port map (
            O => \N__13088\,
            I => \N__13079\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__13085\,
            I => \N__13076\
        );

    \I__3146\ : Sp12to4
    port map (
            O => \N__13082\,
            I => \N__13073\
        );

    \I__3145\ : Span4Mux_v
    port map (
            O => \N__13079\,
            I => \N__13070\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__13076\,
            I => \N__13067\
        );

    \I__3143\ : Odrv12
    port map (
            O => \N__13073\,
            I => \inst_midgetv_core.INSTR_18\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__13070\,
            I => \inst_midgetv_core.INSTR_18\
        );

    \I__3141\ : Odrv4
    port map (
            O => \N__13067\,
            I => \inst_midgetv_core.INSTR_18\
        );

    \I__3140\ : InMux
    port map (
            O => \N__13060\,
            I => \N__13055\
        );

    \I__3139\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13052\
        );

    \I__3138\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13049\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__13055\,
            I => \N__13046\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__13052\,
            I => \N__13041\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__13049\,
            I => \N__13041\
        );

    \I__3134\ : Span12Mux_s10_v
    port map (
            O => \N__13046\,
            I => \N__13038\
        );

    \I__3133\ : Odrv12
    port map (
            O => \N__13041\,
            I => \inst_midgetv_core.INSTR_23\
        );

    \I__3132\ : Odrv12
    port map (
            O => \N__13038\,
            I => \inst_midgetv_core.INSTR_23\
        );

    \I__3131\ : InMux
    port map (
            O => \N__13033\,
            I => \N__13030\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__13030\,
            I => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_3\
        );

    \I__3129\ : InMux
    port map (
            O => \N__13027\,
            I => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_2\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__13024\,
            I => \N__13021\
        );

    \I__3127\ : InMux
    port map (
            O => \N__13021\,
            I => \N__13018\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__13018\,
            I => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_4\
        );

    \I__3125\ : InMux
    port map (
            O => \N__13015\,
            I => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_3\
        );

    \I__3124\ : SRMux
    port map (
            O => \N__13012\,
            I => \N__13005\
        );

    \I__3123\ : SRMux
    port map (
            O => \N__13011\,
            I => \N__13002\
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__13010\,
            I => \N__12999\
        );

    \I__3121\ : SRMux
    port map (
            O => \N__13009\,
            I => \N__12986\
        );

    \I__3120\ : SRMux
    port map (
            O => \N__13008\,
            I => \N__12979\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__13005\,
            I => \N__12975\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__13002\,
            I => \N__12972\
        );

    \I__3117\ : InMux
    port map (
            O => \N__12999\,
            I => \N__12969\
        );

    \I__3116\ : InMux
    port map (
            O => \N__12998\,
            I => \N__12966\
        );

    \I__3115\ : InMux
    port map (
            O => \N__12997\,
            I => \N__12960\
        );

    \I__3114\ : InMux
    port map (
            O => \N__12996\,
            I => \N__12960\
        );

    \I__3113\ : InMux
    port map (
            O => \N__12995\,
            I => \N__12947\
        );

    \I__3112\ : InMux
    port map (
            O => \N__12994\,
            I => \N__12947\
        );

    \I__3111\ : InMux
    port map (
            O => \N__12993\,
            I => \N__12947\
        );

    \I__3110\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12947\
        );

    \I__3109\ : InMux
    port map (
            O => \N__12991\,
            I => \N__12947\
        );

    \I__3108\ : InMux
    port map (
            O => \N__12990\,
            I => \N__12947\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__12989\,
            I => \N__12944\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__12986\,
            I => \N__12941\
        );

    \I__3105\ : SRMux
    port map (
            O => \N__12985\,
            I => \N__12938\
        );

    \I__3104\ : SRMux
    port map (
            O => \N__12984\,
            I => \N__12935\
        );

    \I__3103\ : SRMux
    port map (
            O => \N__12983\,
            I => \N__12932\
        );

    \I__3102\ : SRMux
    port map (
            O => \N__12982\,
            I => \N__12929\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__12979\,
            I => \N__12923\
        );

    \I__3100\ : SRMux
    port map (
            O => \N__12978\,
            I => \N__12920\
        );

    \I__3099\ : Span4Mux_v
    port map (
            O => \N__12975\,
            I => \N__12911\
        );

    \I__3098\ : Span4Mux_h
    port map (
            O => \N__12972\,
            I => \N__12911\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__12969\,
            I => \N__12911\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__12966\,
            I => \N__12911\
        );

    \I__3095\ : SRMux
    port map (
            O => \N__12965\,
            I => \N__12908\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__12960\,
            I => \N__12900\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__12947\,
            I => \N__12900\
        );

    \I__3092\ : InMux
    port map (
            O => \N__12944\,
            I => \N__12897\
        );

    \I__3091\ : Span4Mux_s1_v
    port map (
            O => \N__12941\,
            I => \N__12890\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__12938\,
            I => \N__12890\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__12935\,
            I => \N__12890\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__12932\,
            I => \N__12885\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__12929\,
            I => \N__12885\
        );

    \I__3086\ : SRMux
    port map (
            O => \N__12928\,
            I => \N__12882\
        );

    \I__3085\ : SRMux
    port map (
            O => \N__12927\,
            I => \N__12879\
        );

    \I__3084\ : SRMux
    port map (
            O => \N__12926\,
            I => \N__12876\
        );

    \I__3083\ : Span4Mux_v
    port map (
            O => \N__12923\,
            I => \N__12867\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__12920\,
            I => \N__12867\
        );

    \I__3081\ : Span4Mux_h
    port map (
            O => \N__12911\,
            I => \N__12867\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__12908\,
            I => \N__12867\
        );

    \I__3079\ : SRMux
    port map (
            O => \N__12907\,
            I => \N__12864\
        );

    \I__3078\ : InMux
    port map (
            O => \N__12906\,
            I => \N__12860\
        );

    \I__3077\ : SRMux
    port map (
            O => \N__12905\,
            I => \N__12857\
        );

    \I__3076\ : Span4Mux_h
    port map (
            O => \N__12900\,
            I => \N__12852\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__12897\,
            I => \N__12852\
        );

    \I__3074\ : Span4Mux_v
    port map (
            O => \N__12890\,
            I => \N__12843\
        );

    \I__3073\ : Span4Mux_v
    port map (
            O => \N__12885\,
            I => \N__12843\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__12882\,
            I => \N__12843\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__12879\,
            I => \N__12843\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__12876\,
            I => \N__12836\
        );

    \I__3069\ : Span4Mux_v
    port map (
            O => \N__12867\,
            I => \N__12836\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__12864\,
            I => \N__12836\
        );

    \I__3067\ : SRMux
    port map (
            O => \N__12863\,
            I => \N__12833\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__12860\,
            I => \N__12830\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__12857\,
            I => \N__12827\
        );

    \I__3064\ : Sp12to4
    port map (
            O => \N__12852\,
            I => \N__12824\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__12843\,
            I => \N__12819\
        );

    \I__3062\ : Span4Mux_v
    port map (
            O => \N__12836\,
            I => \N__12819\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__12833\,
            I => \N__12816\
        );

    \I__3060\ : Span4Mux_h
    port map (
            O => \N__12830\,
            I => \N__12813\
        );

    \I__3059\ : Span4Mux_v
    port map (
            O => \N__12827\,
            I => \N__12810\
        );

    \I__3058\ : Span12Mux_v
    port map (
            O => \N__12824\,
            I => \N__12803\
        );

    \I__3057\ : Sp12to4
    port map (
            O => \N__12819\,
            I => \N__12803\
        );

    \I__3056\ : Sp12to4
    port map (
            O => \N__12816\,
            I => \N__12803\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__12813\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3054\ : Odrv4
    port map (
            O => \N__12810\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3053\ : Odrv12
    port map (
            O => \N__12803\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3052\ : InMux
    port map (
            O => \N__12796\,
            I => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_4\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__12793\,
            I => \N__12790\
        );

    \I__3050\ : InMux
    port map (
            O => \N__12790\,
            I => \N__12785\
        );

    \I__3049\ : InMux
    port map (
            O => \N__12789\,
            I => \N__12782\
        );

    \I__3048\ : InMux
    port map (
            O => \N__12788\,
            I => \N__12779\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__12785\,
            I => \N__12776\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__12782\,
            I => \N__12773\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__12779\,
            I => \N__12770\
        );

    \I__3044\ : Span4Mux_v
    port map (
            O => \N__12776\,
            I => \N__12767\
        );

    \I__3043\ : Span4Mux_h
    port map (
            O => \N__12773\,
            I => \N__12764\
        );

    \I__3042\ : Odrv12
    port map (
            O => \N__12770\,
            I => \inst_midgetv_core.lastshift\
        );

    \I__3041\ : Odrv4
    port map (
            O => \N__12767\,
            I => \inst_midgetv_core.lastshift\
        );

    \I__3040\ : Odrv4
    port map (
            O => \N__12764\,
            I => \inst_midgetv_core.lastshift\
        );

    \I__3039\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12754\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__12754\,
            I => \inst_midgetv_core.inst_shiftcounter.genblk1_d_2\
        );

    \I__3037\ : InMux
    port map (
            O => \N__12751\,
            I => \N__12747\
        );

    \I__3036\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12744\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__12747\,
            I => \N__12739\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__12744\,
            I => \N__12739\
        );

    \I__3033\ : Span4Mux_v
    port map (
            O => \N__12739\,
            I => \N__12735\
        );

    \I__3032\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12732\
        );

    \I__3031\ : Span4Mux_h
    port map (
            O => \N__12735\,
            I => \N__12722\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__12732\,
            I => \N__12719\
        );

    \I__3029\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12714\
        );

    \I__3028\ : InMux
    port map (
            O => \N__12730\,
            I => \N__12714\
        );

    \I__3027\ : InMux
    port map (
            O => \N__12729\,
            I => \N__12709\
        );

    \I__3026\ : InMux
    port map (
            O => \N__12728\,
            I => \N__12709\
        );

    \I__3025\ : InMux
    port map (
            O => \N__12727\,
            I => \N__12706\
        );

    \I__3024\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12703\
        );

    \I__3023\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12700\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__12722\,
            I => \N__12697\
        );

    \I__3021\ : Span4Mux_v
    port map (
            O => \N__12719\,
            I => \N__12690\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__12714\,
            I => \N__12690\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__12709\,
            I => \N__12690\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__12706\,
            I => \N__12687\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__12703\,
            I => \N__12682\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__12700\,
            I => \N__12682\
        );

    \I__3015\ : Sp12to4
    port map (
            O => \N__12697\,
            I => \N__12679\
        );

    \I__3014\ : Span4Mux_h
    port map (
            O => \N__12690\,
            I => \N__12674\
        );

    \I__3013\ : Span4Mux_v
    port map (
            O => \N__12687\,
            I => \N__12674\
        );

    \I__3012\ : Span12Mux_v
    port map (
            O => \N__12682\,
            I => \N__12669\
        );

    \I__3011\ : Span12Mux_v
    port map (
            O => \N__12679\,
            I => \N__12669\
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__12674\,
            I => \inst_midgetv_core.B_1\
        );

    \I__3009\ : Odrv12
    port map (
            O => \N__12669\,
            I => \inst_midgetv_core.B_1\
        );

    \I__3008\ : InMux
    port map (
            O => \N__12664\,
            I => \N__12661\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__12661\,
            I => \inst_midgetv_core.inst_shiftcounter.genblk1_d_3\
        );

    \I__3006\ : InMux
    port map (
            O => \N__12658\,
            I => \N__12655\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__12655\,
            I => \N__12652\
        );

    \I__3004\ : Odrv4
    port map (
            O => \N__12652\,
            I => \inst_midgetv_core.bmask_2\
        );

    \I__3003\ : CEMux
    port map (
            O => \N__12649\,
            I => \N__12646\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__12646\,
            I => \N__12642\
        );

    \I__3001\ : CEMux
    port map (
            O => \N__12645\,
            I => \N__12639\
        );

    \I__3000\ : Span4Mux_v
    port map (
            O => \N__12642\,
            I => \N__12634\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__12639\,
            I => \N__12634\
        );

    \I__2998\ : Span4Mux_v
    port map (
            O => \N__12634\,
            I => \N__12631\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__12631\,
            I => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.we\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__12628\,
            I => \N__12625\
        );

    \I__2995\ : InMux
    port map (
            O => \N__12625\,
            I => \N__12622\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__12622\,
            I => \inst_midgetv_core.bmask_3\
        );

    \I__2993\ : CEMux
    port map (
            O => \N__12619\,
            I => \N__12615\
        );

    \I__2992\ : CEMux
    port map (
            O => \N__12618\,
            I => \N__12612\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__12615\,
            I => \N__12607\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__12612\,
            I => \N__12607\
        );

    \I__2989\ : Span4Mux_s3_v
    port map (
            O => \N__12607\,
            I => \N__12604\
        );

    \I__2988\ : Span4Mux_v
    port map (
            O => \N__12604\,
            I => \N__12601\
        );

    \I__2987\ : Span4Mux_v
    port map (
            O => \N__12601\,
            I => \N__12598\
        );

    \I__2986\ : Odrv4
    port map (
            O => \N__12598\,
            I => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.we\
        );

    \I__2985\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12592\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__12592\,
            I => \N__12589\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__12589\,
            I => \inst_midgetv_core.bmask_1\
        );

    \I__2982\ : InMux
    port map (
            O => \N__12586\,
            I => \N__12577\
        );

    \I__2981\ : InMux
    port map (
            O => \N__12585\,
            I => \N__12577\
        );

    \I__2980\ : InMux
    port map (
            O => \N__12584\,
            I => \N__12577\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__12577\,
            I => \N__12573\
        );

    \I__2978\ : InMux
    port map (
            O => \N__12576\,
            I => \N__12570\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__12573\,
            I => \inst_midgetv_core.iwe\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__12570\,
            I => \inst_midgetv_core.iwe\
        );

    \I__2975\ : CEMux
    port map (
            O => \N__12565\,
            I => \N__12562\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__12562\,
            I => \N__12558\
        );

    \I__2973\ : CEMux
    port map (
            O => \N__12561\,
            I => \N__12555\
        );

    \I__2972\ : Span4Mux_v
    port map (
            O => \N__12558\,
            I => \N__12550\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__12555\,
            I => \N__12550\
        );

    \I__2970\ : Span4Mux_h
    port map (
            O => \N__12550\,
            I => \N__12547\
        );

    \I__2969\ : Span4Mux_h
    port map (
            O => \N__12547\,
            I => \N__12544\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__12544\,
            I => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.we\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__12541\,
            I => \N__12536\
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__12540\,
            I => \N__12531\
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__12539\,
            I => \N__12527\
        );

    \I__2964\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12524\
        );

    \I__2963\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12513\
        );

    \I__2962\ : InMux
    port map (
            O => \N__12534\,
            I => \N__12513\
        );

    \I__2961\ : InMux
    port map (
            O => \N__12531\,
            I => \N__12513\
        );

    \I__2960\ : InMux
    port map (
            O => \N__12530\,
            I => \N__12513\
        );

    \I__2959\ : InMux
    port map (
            O => \N__12527\,
            I => \N__12513\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__12524\,
            I => \N__12510\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__12513\,
            I => \N__12507\
        );

    \I__2956\ : Sp12to4
    port map (
            O => \N__12510\,
            I => \N__12502\
        );

    \I__2955\ : Sp12to4
    port map (
            O => \N__12507\,
            I => \N__12502\
        );

    \I__2954\ : Odrv12
    port map (
            O => \N__12502\,
            I => \inst_midgetv_core.s_shift_1\
        );

    \I__2953\ : InMux
    port map (
            O => \N__12499\,
            I => \N__12496\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__12496\,
            I => \N__12489\
        );

    \I__2951\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12486\
        );

    \I__2950\ : InMux
    port map (
            O => \N__12494\,
            I => \N__12483\
        );

    \I__2949\ : InMux
    port map (
            O => \N__12493\,
            I => \N__12480\
        );

    \I__2948\ : InMux
    port map (
            O => \N__12492\,
            I => \N__12474\
        );

    \I__2947\ : Span4Mux_v
    port map (
            O => \N__12489\,
            I => \N__12466\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__12486\,
            I => \N__12466\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__12483\,
            I => \N__12466\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__12480\,
            I => \N__12462\
        );

    \I__2943\ : InMux
    port map (
            O => \N__12479\,
            I => \N__12457\
        );

    \I__2942\ : InMux
    port map (
            O => \N__12478\,
            I => \N__12457\
        );

    \I__2941\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12454\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__12474\,
            I => \N__12451\
        );

    \I__2939\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12448\
        );

    \I__2938\ : Span4Mux_v
    port map (
            O => \N__12466\,
            I => \N__12445\
        );

    \I__2937\ : InMux
    port map (
            O => \N__12465\,
            I => \N__12442\
        );

    \I__2936\ : Span12Mux_v
    port map (
            O => \N__12462\,
            I => \N__12435\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__12457\,
            I => \N__12435\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__12454\,
            I => \N__12435\
        );

    \I__2933\ : Span4Mux_h
    port map (
            O => \N__12451\,
            I => \N__12432\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__12448\,
            I => \N__12429\
        );

    \I__2931\ : Span4Mux_h
    port map (
            O => \N__12445\,
            I => \N__12424\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__12442\,
            I => \N__12424\
        );

    \I__2929\ : Odrv12
    port map (
            O => \N__12435\,
            I => \inst_midgetv_core.B_0\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__12432\,
            I => \inst_midgetv_core.B_0\
        );

    \I__2927\ : Odrv12
    port map (
            O => \N__12429\,
            I => \inst_midgetv_core.B_0\
        );

    \I__2926\ : Odrv4
    port map (
            O => \N__12424\,
            I => \inst_midgetv_core.B_0\
        );

    \I__2925\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12412\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__12412\,
            I => \N__12409\
        );

    \I__2923\ : Span4Mux_h
    port map (
            O => \N__12409\,
            I => \N__12406\
        );

    \I__2922\ : Span4Mux_h
    port map (
            O => \N__12406\,
            I => \N__12403\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__12403\,
            I => \inst_midgetv_core.s_alu_carryin_0\
        );

    \I__2920\ : InMux
    port map (
            O => \N__12400\,
            I => \N__12396\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__12399\,
            I => \N__12393\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__12396\,
            I => \N__12386\
        );

    \I__2917\ : InMux
    port map (
            O => \N__12393\,
            I => \N__12379\
        );

    \I__2916\ : InMux
    port map (
            O => \N__12392\,
            I => \N__12379\
        );

    \I__2915\ : InMux
    port map (
            O => \N__12391\,
            I => \N__12379\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__12390\,
            I => \N__12376\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__12389\,
            I => \N__12372\
        );

    \I__2912\ : Span4Mux_h
    port map (
            O => \N__12386\,
            I => \N__12364\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__12379\,
            I => \N__12361\
        );

    \I__2910\ : InMux
    port map (
            O => \N__12376\,
            I => \N__12352\
        );

    \I__2909\ : InMux
    port map (
            O => \N__12375\,
            I => \N__12352\
        );

    \I__2908\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12352\
        );

    \I__2907\ : InMux
    port map (
            O => \N__12371\,
            I => \N__12352\
        );

    \I__2906\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12343\
        );

    \I__2905\ : InMux
    port map (
            O => \N__12369\,
            I => \N__12343\
        );

    \I__2904\ : InMux
    port map (
            O => \N__12368\,
            I => \N__12343\
        );

    \I__2903\ : InMux
    port map (
            O => \N__12367\,
            I => \N__12343\
        );

    \I__2902\ : Odrv4
    port map (
            O => \N__12364\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_28\
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__12361\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_28\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__12352\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_28\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__12343\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_28\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__12334\,
            I => \N__12331\
        );

    \I__2897\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12328\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__12328\,
            I => \N__12321\
        );

    \I__2895\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12314\
        );

    \I__2894\ : InMux
    port map (
            O => \N__12326\,
            I => \N__12314\
        );

    \I__2893\ : InMux
    port map (
            O => \N__12325\,
            I => \N__12314\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__12324\,
            I => \N__12308\
        );

    \I__2891\ : Span4Mux_v
    port map (
            O => \N__12321\,
            I => \N__12299\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__12314\,
            I => \N__12299\
        );

    \I__2889\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12290\
        );

    \I__2888\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12290\
        );

    \I__2887\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12290\
        );

    \I__2886\ : InMux
    port map (
            O => \N__12308\,
            I => \N__12290\
        );

    \I__2885\ : InMux
    port map (
            O => \N__12307\,
            I => \N__12281\
        );

    \I__2884\ : InMux
    port map (
            O => \N__12306\,
            I => \N__12281\
        );

    \I__2883\ : InMux
    port map (
            O => \N__12305\,
            I => \N__12281\
        );

    \I__2882\ : InMux
    port map (
            O => \N__12304\,
            I => \N__12281\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__12299\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_31\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__12290\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_31\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__12281\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_31\
        );

    \I__2878\ : InMux
    port map (
            O => \N__12274\,
            I => \N__12269\
        );

    \I__2877\ : CascadeMux
    port map (
            O => \N__12273\,
            I => \N__12266\
        );

    \I__2876\ : CascadeMux
    port map (
            O => \N__12272\,
            I => \N__12263\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__12269\,
            I => \N__12258\
        );

    \I__2874\ : InMux
    port map (
            O => \N__12266\,
            I => \N__12251\
        );

    \I__2873\ : InMux
    port map (
            O => \N__12263\,
            I => \N__12251\
        );

    \I__2872\ : InMux
    port map (
            O => \N__12262\,
            I => \N__12251\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__12261\,
            I => \N__12244\
        );

    \I__2870\ : Span4Mux_v
    port map (
            O => \N__12258\,
            I => \N__12236\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__12251\,
            I => \N__12236\
        );

    \I__2868\ : InMux
    port map (
            O => \N__12250\,
            I => \N__12227\
        );

    \I__2867\ : InMux
    port map (
            O => \N__12249\,
            I => \N__12227\
        );

    \I__2866\ : InMux
    port map (
            O => \N__12248\,
            I => \N__12227\
        );

    \I__2865\ : InMux
    port map (
            O => \N__12247\,
            I => \N__12227\
        );

    \I__2864\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12224\
        );

    \I__2863\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12217\
        );

    \I__2862\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12217\
        );

    \I__2861\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12217\
        );

    \I__2860\ : Odrv4
    port map (
            O => \N__12236\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_30\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__12227\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_30\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__12224\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_30\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__12217\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_30\
        );

    \I__2856\ : InMux
    port map (
            O => \N__12208\,
            I => \N__12205\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__12205\,
            I => \N__12194\
        );

    \I__2854\ : InMux
    port map (
            O => \N__12204\,
            I => \N__12187\
        );

    \I__2853\ : InMux
    port map (
            O => \N__12203\,
            I => \N__12187\
        );

    \I__2852\ : InMux
    port map (
            O => \N__12202\,
            I => \N__12187\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__12201\,
            I => \N__12184\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__12200\,
            I => \N__12181\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__12199\,
            I => \N__12177\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__12198\,
            I => \N__12173\
        );

    \I__2847\ : InMux
    port map (
            O => \N__12197\,
            I => \N__12169\
        );

    \I__2846\ : Span4Mux_h
    port map (
            O => \N__12194\,
            I => \N__12166\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__12187\,
            I => \N__12163\
        );

    \I__2844\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12156\
        );

    \I__2843\ : InMux
    port map (
            O => \N__12181\,
            I => \N__12156\
        );

    \I__2842\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12156\
        );

    \I__2841\ : InMux
    port map (
            O => \N__12177\,
            I => \N__12147\
        );

    \I__2840\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12147\
        );

    \I__2839\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12147\
        );

    \I__2838\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12147\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__12169\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_29\
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__12166\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_29\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__12163\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_29\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__12156\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_29\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__12147\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.indir_29\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__12136\,
            I => \N__12133\
        );

    \I__2831\ : InMux
    port map (
            O => \N__12133\,
            I => \N__12130\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__12130\,
            I => \N__12127\
        );

    \I__2829\ : Span4Mux_v
    port map (
            O => \N__12127\,
            I => \N__12124\
        );

    \I__2828\ : Span4Mux_h
    port map (
            O => \N__12124\,
            I => \N__12121\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__12121\,
            I => \inst_midgetv_core.s_alu_carryin_1\
        );

    \I__2826\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12112\
        );

    \I__2825\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12106\
        );

    \I__2824\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12106\
        );

    \I__2823\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12103\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__12112\,
            I => \N__12099\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__12111\,
            I => \N__12096\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__12106\,
            I => \N__12091\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__12103\,
            I => \N__12091\
        );

    \I__2818\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12088\
        );

    \I__2817\ : Span4Mux_h
    port map (
            O => \N__12099\,
            I => \N__12085\
        );

    \I__2816\ : InMux
    port map (
            O => \N__12096\,
            I => \N__12082\
        );

    \I__2815\ : Span4Mux_v
    port map (
            O => \N__12091\,
            I => \N__12079\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__12088\,
            I => \inst_midgetv_core.sa24\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__12085\,
            I => \inst_midgetv_core.sa24\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__12082\,
            I => \inst_midgetv_core.sa24\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__12079\,
            I => \inst_midgetv_core.sa24\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__12070\,
            I => \N__12065\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__12069\,
            I => \N__12062\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__12068\,
            I => \N__12059\
        );

    \I__2807\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12053\
        );

    \I__2806\ : InMux
    port map (
            O => \N__12062\,
            I => \N__12053\
        );

    \I__2805\ : InMux
    port map (
            O => \N__12059\,
            I => \N__12050\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__12058\,
            I => \N__12047\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__12053\,
            I => \N__12044\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__12050\,
            I => \N__12041\
        );

    \I__2801\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12038\
        );

    \I__2800\ : Span4Mux_v
    port map (
            O => \N__12044\,
            I => \N__12035\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__12041\,
            I => \inst_midgetv_core.inst_progressctrl.blka_usedefault\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__12038\,
            I => \inst_midgetv_core.inst_progressctrl.blka_usedefault\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__12035\,
            I => \inst_midgetv_core.inst_progressctrl.blka_usedefault\
        );

    \I__2796\ : CEMux
    port map (
            O => \N__12028\,
            I => \N__12023\
        );

    \I__2795\ : CEMux
    port map (
            O => \N__12027\,
            I => \N__12020\
        );

    \I__2794\ : CEMux
    port map (
            O => \N__12026\,
            I => \N__12017\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__12023\,
            I => \N__12014\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__12020\,
            I => \N__12011\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__12017\,
            I => \N__12008\
        );

    \I__2790\ : Span4Mux_v
    port map (
            O => \N__12014\,
            I => \N__12003\
        );

    \I__2789\ : Span4Mux_h
    port map (
            O => \N__12011\,
            I => \N__12003\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__12008\,
            I => \inst_midgetv_core.inst_progressctrl.blka_en\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__12003\,
            I => \inst_midgetv_core.inst_progressctrl.blka_en\
        );

    \I__2786\ : InMux
    port map (
            O => \N__11998\,
            I => \N__11995\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__11995\,
            I => \inst_midgetv_core.inst_shiftcounter.genblk1_d_0\
        );

    \I__2784\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11989\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__11989\,
            I => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_1\
        );

    \I__2782\ : InMux
    port map (
            O => \N__11986\,
            I => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_0\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__11983\,
            I => \N__11980\
        );

    \I__2780\ : InMux
    port map (
            O => \N__11980\,
            I => \N__11977\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__11977\,
            I => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_2\
        );

    \I__2778\ : InMux
    port map (
            O => \N__11974\,
            I => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_1\
        );

    \I__2777\ : SRMux
    port map (
            O => \N__11971\,
            I => \N__11968\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__11968\,
            I => \N__11965\
        );

    \I__2775\ : Span4Mux_h
    port map (
            O => \N__11965\,
            I => \N__11961\
        );

    \I__2774\ : InMux
    port map (
            O => \N__11964\,
            I => \N__11958\
        );

    \I__2773\ : Span4Mux_v
    port map (
            O => \N__11961\,
            I => \N__11953\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__11958\,
            I => \N__11950\
        );

    \I__2771\ : InMux
    port map (
            O => \N__11957\,
            I => \N__11945\
        );

    \I__2770\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11945\
        );

    \I__2769\ : Span4Mux_h
    port map (
            O => \N__11953\,
            I => \N__11939\
        );

    \I__2768\ : Span4Mux_h
    port map (
            O => \N__11950\,
            I => \N__11939\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__11945\,
            I => \N__11936\
        );

    \I__2766\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11933\
        );

    \I__2765\ : Odrv4
    port map (
            O => \N__11939\,
            I => \inst_midgetv_core.buserror\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__11936\,
            I => \inst_midgetv_core.buserror\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__11933\,
            I => \inst_midgetv_core.buserror\
        );

    \I__2762\ : CEMux
    port map (
            O => \N__11926\,
            I => \N__11923\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__11923\,
            I => \N__11920\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__11920\,
            I => \N__11916\
        );

    \I__2759\ : CEMux
    port map (
            O => \N__11919\,
            I => \N__11913\
        );

    \I__2758\ : Sp12to4
    port map (
            O => \N__11916\,
            I => \N__11908\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__11913\,
            I => \N__11908\
        );

    \I__2756\ : Odrv12
    port map (
            O => \N__11908\,
            I => \CONSTANT_ZERO_NET\
        );

    \I__2755\ : InMux
    port map (
            O => \N__11905\,
            I => \N__11902\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__11902\,
            I => \N__11898\
        );

    \I__2753\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11895\
        );

    \I__2752\ : Span4Mux_h
    port map (
            O => \N__11898\,
            I => \N__11890\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__11895\,
            I => \N__11890\
        );

    \I__2750\ : Odrv4
    port map (
            O => \N__11890\,
            I => \inst_midgetv_core.sa15\
        );

    \I__2749\ : InMux
    port map (
            O => \N__11887\,
            I => \N__11883\
        );

    \I__2748\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11880\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__11883\,
            I => \inst_midgetv_core.sa32\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__11880\,
            I => \inst_midgetv_core.sa32\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__11875\,
            I => \N__11872\
        );

    \I__2744\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11869\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__11869\,
            I => \N__11865\
        );

    \I__2742\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11862\
        );

    \I__2741\ : Odrv12
    port map (
            O => \N__11865\,
            I => \inst_midgetv_core.inst_ucodepc.maybranch_N_253\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__11862\,
            I => \inst_midgetv_core.inst_ucodepc.maybranch_N_253\
        );

    \I__2739\ : InMux
    port map (
            O => \N__11857\,
            I => \N__11854\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__11854\,
            I => \N__11850\
        );

    \I__2737\ : InMux
    port map (
            O => \N__11853\,
            I => \N__11847\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__11850\,
            I => \N__11843\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__11847\,
            I => \N__11840\
        );

    \I__2734\ : InMux
    port map (
            O => \N__11846\,
            I => \N__11837\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__11843\,
            I => \inst_midgetv_core.sa30\
        );

    \I__2732\ : Odrv12
    port map (
            O => \N__11840\,
            I => \inst_midgetv_core.sa30\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__11837\,
            I => \inst_midgetv_core.sa30\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__11830\,
            I => \N__11827\
        );

    \I__2729\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11824\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__11824\,
            I => \N__11820\
        );

    \I__2727\ : InMux
    port map (
            O => \N__11823\,
            I => \N__11817\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__11820\,
            I => \inst_midgetv_core.sa37\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__11817\,
            I => \inst_midgetv_core.sa37\
        );

    \I__2724\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11806\
        );

    \I__2723\ : InMux
    port map (
            O => \N__11811\,
            I => \N__11806\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__11806\,
            I => \inst_midgetv_core.sa25\
        );

    \I__2721\ : InMux
    port map (
            O => \N__11803\,
            I => \N__11796\
        );

    \I__2720\ : InMux
    port map (
            O => \N__11802\,
            I => \N__11796\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11791\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__11796\,
            I => \N__11788\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11785\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11794\,
            I => \N__11782\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__11791\,
            I => \N__11778\
        );

    \I__2714\ : Span4Mux_v
    port map (
            O => \N__11788\,
            I => \N__11771\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__11785\,
            I => \N__11771\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__11782\,
            I => \N__11771\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__11781\,
            I => \N__11766\
        );

    \I__2710\ : Span4Mux_h
    port map (
            O => \N__11778\,
            I => \N__11763\
        );

    \I__2709\ : Span4Mux_v
    port map (
            O => \N__11771\,
            I => \N__11760\
        );

    \I__2708\ : InMux
    port map (
            O => \N__11770\,
            I => \N__11757\
        );

    \I__2707\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11752\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11766\,
            I => \N__11752\
        );

    \I__2705\ : Odrv4
    port map (
            O => \N__11763\,
            I => \ADR_O_3\
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__11760\,
            I => \ADR_O_3\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11757\,
            I => \ADR_O_3\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__11752\,
            I => \ADR_O_3\
        );

    \I__2701\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11740\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__11740\,
            I => \inst_midgetv_core.inst_wai.genblk1_preWai1\
        );

    \I__2699\ : InMux
    port map (
            O => \N__11737\,
            I => \N__11733\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__11736\,
            I => \N__11730\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__11733\,
            I => \N__11727\
        );

    \I__2696\ : InMux
    port map (
            O => \N__11730\,
            I => \N__11724\
        );

    \I__2695\ : Span4Mux_h
    port map (
            O => \N__11727\,
            I => \N__11717\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__11724\,
            I => \N__11717\
        );

    \I__2693\ : InMux
    port map (
            O => \N__11723\,
            I => \N__11712\
        );

    \I__2692\ : InMux
    port map (
            O => \N__11722\,
            I => \N__11712\
        );

    \I__2691\ : Odrv4
    port map (
            O => \N__11717\,
            I => \inst_midgetv_core.ADR_O_11\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__11712\,
            I => \inst_midgetv_core.ADR_O_11\
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__11707\,
            I => \N__11704\
        );

    \I__2688\ : CascadeBuf
    port map (
            O => \N__11704\,
            I => \N__11701\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__11701\,
            I => \N__11698\
        );

    \I__2686\ : CascadeBuf
    port map (
            O => \N__11698\,
            I => \N__11695\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__11695\,
            I => \N__11692\
        );

    \I__2684\ : CascadeBuf
    port map (
            O => \N__11692\,
            I => \N__11689\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__11689\,
            I => \N__11686\
        );

    \I__2682\ : CascadeBuf
    port map (
            O => \N__11686\,
            I => \N__11683\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__11683\,
            I => \N__11680\
        );

    \I__2680\ : CascadeBuf
    port map (
            O => \N__11680\,
            I => \N__11677\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__11677\,
            I => \N__11674\
        );

    \I__2678\ : CascadeBuf
    port map (
            O => \N__11674\,
            I => \N__11671\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__11671\,
            I => \N__11668\
        );

    \I__2676\ : CascadeBuf
    port map (
            O => \N__11668\,
            I => \N__11665\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__11665\,
            I => \N__11662\
        );

    \I__2674\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11659\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__11659\,
            I => \N__11656\
        );

    \I__2672\ : Span12Mux_s8_h
    port map (
            O => \N__11656\,
            I => \N__11653\
        );

    \I__2671\ : Odrv12
    port map (
            O => \N__11653\,
            I => \inst_midgetv_core.Wai_9\
        );

    \I__2670\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11647\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__11647\,
            I => \N__11644\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__11644\,
            I => \SEL_O_3\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11641\,
            I => \N__11638\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__11638\,
            I => \N__11634\
        );

    \I__2665\ : InMux
    port map (
            O => \N__11637\,
            I => \N__11631\
        );

    \I__2664\ : Span4Mux_h
    port map (
            O => \N__11634\,
            I => \N__11628\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11631\,
            I => \N__11625\
        );

    \I__2662\ : Span4Mux_v
    port map (
            O => \N__11628\,
            I => \N__11622\
        );

    \I__2661\ : Span12Mux_h
    port map (
            O => \N__11625\,
            I => \N__11619\
        );

    \I__2660\ : Span4Mux_v
    port map (
            O => \N__11622\,
            I => \N__11616\
        );

    \I__2659\ : Odrv12
    port map (
            O => \N__11619\,
            I => \DAT_O_31\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__11616\,
            I => \DAT_O_31\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__11611\,
            I => \N__11607\
        );

    \I__2656\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11603\
        );

    \I__2655\ : InMux
    port map (
            O => \N__11607\,
            I => \N__11598\
        );

    \I__2654\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11598\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__11603\,
            I => bluesource_is_uart
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__11598\,
            I => bluesource_is_uart
        );

    \I__2651\ : CEMux
    port map (
            O => \N__11593\,
            I => \N__11590\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__11590\,
            I => \N__11587\
        );

    \I__2649\ : Sp12to4
    port map (
            O => \N__11587\,
            I => \N__11584\
        );

    \I__2648\ : Odrv12
    port map (
            O => \N__11584\,
            I => \i_LEDs.n2766\
        );

    \I__2647\ : CEMux
    port map (
            O => \N__11581\,
            I => \N__11578\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11578\,
            I => \N__11575\
        );

    \I__2645\ : IoSpan4Mux
    port map (
            O => \N__11575\,
            I => \N__11572\
        );

    \I__2644\ : Span4Mux_s1_v
    port map (
            O => \N__11572\,
            I => \N__11569\
        );

    \I__2643\ : Sp12to4
    port map (
            O => \N__11569\,
            I => \N__11566\
        );

    \I__2642\ : Span12Mux_s9_v
    port map (
            O => \N__11566\,
            I => \N__11563\
        );

    \I__2641\ : Odrv12
    port map (
            O => \N__11563\,
            I => \i_BBUART.usartTX_N_2\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11560\,
            I => \N__11555\
        );

    \I__2639\ : InMux
    port map (
            O => \N__11559\,
            I => \N__11550\
        );

    \I__2638\ : InMux
    port map (
            O => \N__11558\,
            I => \N__11550\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__11555\,
            I => \N__11547\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__11550\,
            I => \N__11542\
        );

    \I__2635\ : Span4Mux_h
    port map (
            O => \N__11547\,
            I => \N__11542\
        );

    \I__2634\ : Span4Mux_v
    port map (
            O => \N__11542\,
            I => \N__11539\
        );

    \I__2633\ : Odrv4
    port map (
            O => \N__11539\,
            I => \WE_O\
        );

    \I__2632\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11529\
        );

    \I__2631\ : InMux
    port map (
            O => \N__11535\,
            I => \N__11529\
        );

    \I__2630\ : InMux
    port map (
            O => \N__11534\,
            I => \N__11525\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__11529\,
            I => \N__11522\
        );

    \I__2628\ : InMux
    port map (
            O => \N__11528\,
            I => \N__11519\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__11525\,
            I => \N__11516\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__11522\,
            I => \N__11511\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__11519\,
            I => \N__11511\
        );

    \I__2624\ : Span4Mux_h
    port map (
            O => \N__11516\,
            I => \N__11503\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__11511\,
            I => \N__11503\
        );

    \I__2622\ : InMux
    port map (
            O => \N__11510\,
            I => \N__11500\
        );

    \I__2621\ : InMux
    port map (
            O => \N__11509\,
            I => \N__11495\
        );

    \I__2620\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11495\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__11503\,
            I => \ADR_O_2\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__11500\,
            I => \ADR_O_2\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__11495\,
            I => \ADR_O_2\
        );

    \I__2616\ : CEMux
    port map (
            O => \N__11488\,
            I => \N__11485\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__11485\,
            I => \N__11481\
        );

    \I__2614\ : CEMux
    port map (
            O => \N__11484\,
            I => \N__11478\
        );

    \I__2613\ : IoSpan4Mux
    port map (
            O => \N__11481\,
            I => \N__11475\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__11478\,
            I => \N__11472\
        );

    \I__2611\ : Span4Mux_s3_v
    port map (
            O => \N__11475\,
            I => \N__11465\
        );

    \I__2610\ : Span4Mux_s3_v
    port map (
            O => \N__11472\,
            I => \N__11465\
        );

    \I__2609\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11460\
        );

    \I__2608\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11460\
        );

    \I__2607\ : Span4Mux_v
    port map (
            O => \N__11465\,
            I => \N__11457\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__11460\,
            I => \N__11454\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__11457\,
            I => \LED1_N_4\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__11454\,
            I => \LED1_N_4\
        );

    \I__2603\ : InMux
    port map (
            O => \N__11449\,
            I => \N__11446\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__11446\,
            I => \inst_midgetv_core.inst_progressctrl.n4_adj_311\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__11443\,
            I => \N__11440\
        );

    \I__2600\ : InMux
    port map (
            O => \N__11440\,
            I => \N__11437\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__11437\,
            I => n2345
        );

    \I__2598\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11430\
        );

    \I__2597\ : InMux
    port map (
            O => \N__11433\,
            I => \N__11427\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__11430\,
            I => \N__11422\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__11427\,
            I => \N__11419\
        );

    \I__2594\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11412\
        );

    \I__2593\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11412\
        );

    \I__2592\ : Sp12to4
    port map (
            O => \N__11422\,
            I => \N__11409\
        );

    \I__2591\ : Span4Mux_h
    port map (
            O => \N__11419\,
            I => \N__11406\
        );

    \I__2590\ : InMux
    port map (
            O => \N__11418\,
            I => \N__11403\
        );

    \I__2589\ : InMux
    port map (
            O => \N__11417\,
            I => \N__11400\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__11412\,
            I => \N__11395\
        );

    \I__2587\ : Span12Mux_s9_v
    port map (
            O => \N__11409\,
            I => \N__11395\
        );

    \I__2586\ : Span4Mux_h
    port map (
            O => \N__11406\,
            I => \N__11392\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__11403\,
            I => \N__11389\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__11400\,
            I => \inst_midgetv_core.B_31\
        );

    \I__2583\ : Odrv12
    port map (
            O => \N__11395\,
            I => \inst_midgetv_core.B_31\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__11392\,
            I => \inst_midgetv_core.B_31\
        );

    \I__2581\ : Odrv12
    port map (
            O => \N__11389\,
            I => \inst_midgetv_core.B_31\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__11380\,
            I => \N__11377\
        );

    \I__2579\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11374\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__11374\,
            I => \N__11370\
        );

    \I__2577\ : InMux
    port map (
            O => \N__11373\,
            I => \N__11367\
        );

    \I__2576\ : Span4Mux_h
    port map (
            O => \N__11370\,
            I => \N__11362\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__11367\,
            I => \N__11362\
        );

    \I__2574\ : Span4Mux_v
    port map (
            O => \N__11362\,
            I => \N__11359\
        );

    \I__2573\ : Span4Mux_v
    port map (
            O => \N__11359\,
            I => \N__11356\
        );

    \I__2572\ : Odrv4
    port map (
            O => \N__11356\,
            I => \inst_midgetv_core.sa42\
        );

    \I__2571\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11349\
        );

    \I__2570\ : InMux
    port map (
            O => \N__11352\,
            I => \N__11346\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__11349\,
            I => \N__11342\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__11346\,
            I => \N__11339\
        );

    \I__2567\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11336\
        );

    \I__2566\ : Span4Mux_h
    port map (
            O => \N__11342\,
            I => \N__11329\
        );

    \I__2565\ : Span4Mux_h
    port map (
            O => \N__11339\,
            I => \N__11329\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__11336\,
            I => \N__11329\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__11329\,
            I => \N__11326\
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__11326\,
            I => \inst_midgetv_core.inst_progressctrl.badalignment\
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__11323\,
            I => \N__11316\
        );

    \I__2560\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11312\
        );

    \I__2559\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11309\
        );

    \I__2558\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11304\
        );

    \I__2557\ : InMux
    port map (
            O => \N__11319\,
            I => \N__11304\
        );

    \I__2556\ : InMux
    port map (
            O => \N__11316\,
            I => \N__11301\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__11315\,
            I => \N__11297\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__11312\,
            I => \N__11294\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__11309\,
            I => \N__11291\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__11304\,
            I => \N__11288\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__11301\,
            I => \N__11285\
        );

    \I__2550\ : InMux
    port map (
            O => \N__11300\,
            I => \N__11280\
        );

    \I__2549\ : InMux
    port map (
            O => \N__11297\,
            I => \N__11280\
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__11294\,
            I => \inst_midgetv_core.INSTR_6\
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__11291\,
            I => \inst_midgetv_core.INSTR_6\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__11288\,
            I => \inst_midgetv_core.INSTR_6\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__11285\,
            I => \inst_midgetv_core.INSTR_6\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__11280\,
            I => \inst_midgetv_core.INSTR_6\
        );

    \I__2543\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11263\
        );

    \I__2542\ : InMux
    port map (
            O => \N__11268\,
            I => \N__11260\
        );

    \I__2541\ : InMux
    port map (
            O => \N__11267\,
            I => \N__11257\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__11266\,
            I => \N__11253\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__11263\,
            I => \N__11249\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__11260\,
            I => \N__11246\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__11257\,
            I => \N__11238\
        );

    \I__2536\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11231\
        );

    \I__2535\ : InMux
    port map (
            O => \N__11253\,
            I => \N__11231\
        );

    \I__2534\ : InMux
    port map (
            O => \N__11252\,
            I => \N__11231\
        );

    \I__2533\ : Span4Mux_v
    port map (
            O => \N__11249\,
            I => \N__11226\
        );

    \I__2532\ : Span4Mux_v
    port map (
            O => \N__11246\,
            I => \N__11226\
        );

    \I__2531\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11219\
        );

    \I__2530\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11219\
        );

    \I__2529\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11219\
        );

    \I__2528\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11214\
        );

    \I__2527\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11214\
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__11238\,
            I => \inst_midgetv_core.INSTR_2\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__11231\,
            I => \inst_midgetv_core.INSTR_2\
        );

    \I__2524\ : Odrv4
    port map (
            O => \N__11226\,
            I => \inst_midgetv_core.INSTR_2\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__11219\,
            I => \inst_midgetv_core.INSTR_2\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__11214\,
            I => \inst_midgetv_core.INSTR_2\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__11203\,
            I => \N__11199\
        );

    \I__2520\ : InMux
    port map (
            O => \N__11202\,
            I => \N__11194\
        );

    \I__2519\ : InMux
    port map (
            O => \N__11199\,
            I => \N__11191\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__11198\,
            I => \N__11184\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__11197\,
            I => \N__11180\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__11194\,
            I => \N__11176\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__11191\,
            I => \N__11173\
        );

    \I__2514\ : InMux
    port map (
            O => \N__11190\,
            I => \N__11170\
        );

    \I__2513\ : InMux
    port map (
            O => \N__11189\,
            I => \N__11147\
        );

    \I__2512\ : InMux
    port map (
            O => \N__11188\,
            I => \N__11147\
        );

    \I__2511\ : InMux
    port map (
            O => \N__11187\,
            I => \N__11147\
        );

    \I__2510\ : InMux
    port map (
            O => \N__11184\,
            I => \N__11147\
        );

    \I__2509\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11147\
        );

    \I__2508\ : InMux
    port map (
            O => \N__11180\,
            I => \N__11147\
        );

    \I__2507\ : InMux
    port map (
            O => \N__11179\,
            I => \N__11147\
        );

    \I__2506\ : Span4Mux_v
    port map (
            O => \N__11176\,
            I => \N__11144\
        );

    \I__2505\ : Span4Mux_h
    port map (
            O => \N__11173\,
            I => \N__11139\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__11170\,
            I => \N__11139\
        );

    \I__2503\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11128\
        );

    \I__2502\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11128\
        );

    \I__2501\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11128\
        );

    \I__2500\ : InMux
    port map (
            O => \N__11166\,
            I => \N__11128\
        );

    \I__2499\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11128\
        );

    \I__2498\ : InMux
    port map (
            O => \N__11164\,
            I => \N__11121\
        );

    \I__2497\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11121\
        );

    \I__2496\ : InMux
    port map (
            O => \N__11162\,
            I => \N__11121\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__11147\,
            I => \inst_midgetv_core.s_cyclecnt_0\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__11144\,
            I => \inst_midgetv_core.s_cyclecnt_0\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__11139\,
            I => \inst_midgetv_core.s_cyclecnt_0\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__11128\,
            I => \inst_midgetv_core.s_cyclecnt_0\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__11121\,
            I => \inst_midgetv_core.s_cyclecnt_0\
        );

    \I__2490\ : InMux
    port map (
            O => \N__11110\,
            I => \N__11098\
        );

    \I__2489\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11098\
        );

    \I__2488\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11098\
        );

    \I__2487\ : InMux
    port map (
            O => \N__11107\,
            I => \N__11095\
        );

    \I__2486\ : InMux
    port map (
            O => \N__11106\,
            I => \N__11092\
        );

    \I__2485\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11089\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__11098\,
            I => \N__11086\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__11095\,
            I => \N__11078\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__11092\,
            I => \N__11075\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__11089\,
            I => \N__11072\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__11086\,
            I => \N__11069\
        );

    \I__2479\ : InMux
    port map (
            O => \N__11085\,
            I => \N__11066\
        );

    \I__2478\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11059\
        );

    \I__2477\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11059\
        );

    \I__2476\ : InMux
    port map (
            O => \N__11082\,
            I => \N__11059\
        );

    \I__2475\ : InMux
    port map (
            O => \N__11081\,
            I => \N__11056\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__11078\,
            I => \inst_midgetv_core.INSTR_4\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__11075\,
            I => \inst_midgetv_core.INSTR_4\
        );

    \I__2472\ : Odrv4
    port map (
            O => \N__11072\,
            I => \inst_midgetv_core.INSTR_4\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__11069\,
            I => \inst_midgetv_core.INSTR_4\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__11066\,
            I => \inst_midgetv_core.INSTR_4\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__11059\,
            I => \inst_midgetv_core.INSTR_4\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__11056\,
            I => \inst_midgetv_core.INSTR_4\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__11041\,
            I => \N__11038\
        );

    \I__2466\ : InMux
    port map (
            O => \N__11038\,
            I => \N__11034\
        );

    \I__2465\ : InMux
    port map (
            O => \N__11037\,
            I => \N__11030\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__11034\,
            I => \N__11027\
        );

    \I__2463\ : InMux
    port map (
            O => \N__11033\,
            I => \N__11024\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__11030\,
            I => \N__11021\
        );

    \I__2461\ : Span4Mux_h
    port map (
            O => \N__11027\,
            I => \N__11016\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__11024\,
            I => \N__11016\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__11021\,
            I => \inst_midgetv_core.INSTR_8\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__11016\,
            I => \inst_midgetv_core.INSTR_8\
        );

    \I__2457\ : InMux
    port map (
            O => \N__11011\,
            I => \N__11008\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__11008\,
            I => \N__11005\
        );

    \I__2455\ : Span4Mux_h
    port map (
            O => \N__11005\,
            I => \N__11002\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__11002\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm1a\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10999\,
            I => \N__10987\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10987\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10987\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10987\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10987\,
            I => \N__10977\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__10986\,
            I => \N__10974\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__10985\,
            I => \N__10971\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__10984\,
            I => \N__10968\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__10983\,
            I => \N__10965\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__10982\,
            I => \N__10961\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__10981\,
            I => \N__10957\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10950\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__10977\,
            I => \N__10947\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10944\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10971\,
            I => \N__10939\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10968\,
            I => \N__10939\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10932\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10932\
        );

    \I__2435\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10932\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10919\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10957\,
            I => \N__10919\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10919\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10919\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10919\
        );

    \I__2429\ : InMux
    port map (
            O => \N__10953\,
            I => \N__10919\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10950\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09\
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__10947\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__10944\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10939\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10932\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__10919\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10890\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10890\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10890\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10903\,
            I => \N__10890\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__10902\,
            I => \N__10881\
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__10901\,
            I => \N__10877\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10900\,
            I => \N__10874\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10899\,
            I => \N__10871\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__10890\,
            I => \N__10868\
        );

    \I__2413\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10857\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10888\,
            I => \N__10857\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10857\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10857\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10857\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10848\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10848\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10848\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10848\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10874\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa07\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10871\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa07\
        );

    \I__2402\ : Odrv12
    port map (
            O => \N__10868\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa07\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10857\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa07\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10848\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa07\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__10837\,
            I => \N__10833\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__10836\,
            I => \N__10824\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10819\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__10832\,
            I => \N__10816\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__10831\,
            I => \N__10812\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__10830\,
            I => \N__10809\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10796\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10796\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10796\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10796\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10796\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10796\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10819\,
            I => \N__10793\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10790\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10815\,
            I => \N__10783\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10783\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10783\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__10796\,
            I => \N__10780\
        );

    \I__2381\ : Span4Mux_h
    port map (
            O => \N__10793\,
            I => \N__10775\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__10790\,
            I => \N__10775\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10783\,
            I => \N__10770\
        );

    \I__2378\ : Span4Mux_h
    port map (
            O => \N__10780\,
            I => \N__10770\
        );

    \I__2377\ : Span4Mux_h
    port map (
            O => \N__10775\,
            I => \N__10767\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__10770\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa08\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__10767\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa08\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__10762\,
            I => \N__10759\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10759\,
            I => \N__10755\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10758\,
            I => \N__10752\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10755\,
            I => \N__10749\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10752\,
            I => \N__10746\
        );

    \I__2369\ : Span4Mux_v
    port map (
            O => \N__10749\,
            I => \N__10743\
        );

    \I__2368\ : Span4Mux_v
    port map (
            O => \N__10746\,
            I => \N__10737\
        );

    \I__2367\ : Span4Mux_h
    port map (
            O => \N__10743\,
            I => \N__10737\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10742\,
            I => \N__10734\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__10737\,
            I => \inst_midgetv_core.INSTR_10\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__10734\,
            I => \inst_midgetv_core.INSTR_10\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10726\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10726\,
            I => \N__10723\
        );

    \I__2361\ : Span4Mux_v
    port map (
            O => \N__10723\,
            I => \N__10720\
        );

    \I__2360\ : Odrv4
    port map (
            O => \N__10720\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm3a\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10717\,
            I => \N__10714\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__10714\,
            I => \inst_midgetv_core.bmask_0\
        );

    \I__2357\ : CascadeMux
    port map (
            O => \N__10711\,
            I => \N__10708\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10708\,
            I => \N__10705\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__10705\,
            I => \N__10701\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10704\,
            I => \N__10698\
        );

    \I__2353\ : Span4Mux_h
    port map (
            O => \N__10701\,
            I => \N__10695\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__10698\,
            I => \N__10692\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__10695\,
            I => \inst_midgetv_core.rlastshift\
        );

    \I__2350\ : Odrv12
    port map (
            O => \N__10692\,
            I => \inst_midgetv_core.rlastshift\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__10687\,
            I => \N__10683\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10680\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10677\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10680\,
            I => \N__10672\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10677\,
            I => \N__10672\
        );

    \I__2344\ : Span4Mux_v
    port map (
            O => \N__10672\,
            I => \N__10669\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__10669\,
            I => \inst_midgetv_core.sa41\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10663\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__10663\,
            I => \N__10657\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10662\,
            I => \N__10654\
        );

    \I__2339\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10651\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__10660\,
            I => \N__10647\
        );

    \I__2337\ : Span4Mux_v
    port map (
            O => \N__10657\,
            I => \N__10642\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__10654\,
            I => \N__10637\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10651\,
            I => \N__10637\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10650\,
            I => \N__10634\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10631\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10646\,
            I => \N__10626\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10645\,
            I => \N__10626\
        );

    \I__2330\ : Span4Mux_h
    port map (
            O => \N__10642\,
            I => \N__10618\
        );

    \I__2329\ : Span4Mux_v
    port map (
            O => \N__10637\,
            I => \N__10618\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10634\,
            I => \N__10618\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10631\,
            I => \N__10613\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__10626\,
            I => \N__10613\
        );

    \I__2325\ : InMux
    port map (
            O => \N__10625\,
            I => \N__10610\
        );

    \I__2324\ : Span4Mux_h
    port map (
            O => \N__10618\,
            I => \N__10607\
        );

    \I__2323\ : Span4Mux_v
    port map (
            O => \N__10613\,
            I => \N__10604\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__10610\,
            I => corerunning
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__10607\,
            I => corerunning
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__10604\,
            I => corerunning
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__10597\,
            I => \inst_midgetv_core.inst_progressctrl.blka_cmb_bsel_3_cascade_\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10590\
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__10593\,
            I => \N__10587\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__10590\,
            I => \N__10584\
        );

    \I__2315\ : InMux
    port map (
            O => \N__10587\,
            I => \N__10581\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__10584\,
            I => \N__10576\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__10581\,
            I => \N__10576\
        );

    \I__2312\ : Span4Mux_h
    port map (
            O => \N__10576\,
            I => \N__10573\
        );

    \I__2311\ : Span4Mux_v
    port map (
            O => \N__10573\,
            I => \N__10570\
        );

    \I__2310\ : Span4Mux_v
    port map (
            O => \N__10570\,
            I => \N__10567\
        );

    \I__2309\ : Sp12to4
    port map (
            O => \N__10567\,
            I => \N__10564\
        );

    \I__2308\ : Odrv12
    port map (
            O => \N__10564\,
            I => \meta_usartRX\
        );

    \I__2307\ : InMux
    port map (
            O => \N__10561\,
            I => \N__10558\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__10558\,
            I => \N__10554\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10551\
        );

    \I__2304\ : Span4Mux_h
    port map (
            O => \N__10554\,
            I => \N__10548\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__10551\,
            I => \N__10545\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__10548\,
            I => \DAT_O_2\
        );

    \I__2301\ : Odrv12
    port map (
            O => \N__10545\,
            I => \DAT_O_2\
        );

    \I__2300\ : IoInMux
    port map (
            O => \N__10540\,
            I => \N__10537\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__10537\,
            I => \N__10534\
        );

    \I__2298\ : Span4Mux_s0_v
    port map (
            O => \N__10534\,
            I => \N__10531\
        );

    \I__2297\ : Span4Mux_v
    port map (
            O => \N__10531\,
            I => \N__10528\
        );

    \I__2296\ : Span4Mux_v
    port map (
            O => \N__10528\,
            I => \N__10525\
        );

    \I__2295\ : Span4Mux_v
    port map (
            O => \N__10525\,
            I => \N__10522\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__10522\,
            I => \LED3_c\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__10519\,
            I => \N__10516\
        );

    \I__2292\ : CascadeBuf
    port map (
            O => \N__10516\,
            I => \N__10513\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__10513\,
            I => \N__10510\
        );

    \I__2290\ : CascadeBuf
    port map (
            O => \N__10510\,
            I => \N__10507\
        );

    \I__2289\ : CascadeMux
    port map (
            O => \N__10507\,
            I => \N__10504\
        );

    \I__2288\ : CascadeBuf
    port map (
            O => \N__10504\,
            I => \N__10501\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__10501\,
            I => \N__10498\
        );

    \I__2286\ : CascadeBuf
    port map (
            O => \N__10498\,
            I => \N__10495\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__10495\,
            I => \N__10492\
        );

    \I__2284\ : CascadeBuf
    port map (
            O => \N__10492\,
            I => \N__10489\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__10489\,
            I => \N__10486\
        );

    \I__2282\ : CascadeBuf
    port map (
            O => \N__10486\,
            I => \N__10483\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__10483\,
            I => \N__10480\
        );

    \I__2280\ : CascadeBuf
    port map (
            O => \N__10480\,
            I => \N__10477\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__10477\,
            I => \N__10474\
        );

    \I__2278\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10471\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__10471\,
            I => \N__10468\
        );

    \I__2276\ : Span4Mux_s3_v
    port map (
            O => \N__10468\,
            I => \N__10465\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__10465\,
            I => \N__10462\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__10462\,
            I => \N__10459\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__10459\,
            I => \N__10456\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__10456\,
            I => \inst_midgetv_core.Wai_1\
        );

    \I__2271\ : InMux
    port map (
            O => \N__10453\,
            I => \N__10450\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10450\,
            I => \N__10444\
        );

    \I__2269\ : InMux
    port map (
            O => \N__10449\,
            I => \N__10441\
        );

    \I__2268\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10438\
        );

    \I__2267\ : InMux
    port map (
            O => \N__10447\,
            I => \N__10435\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__10444\,
            I => \inst_midgetv_core.ADR_O_4\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__10441\,
            I => \inst_midgetv_core.ADR_O_4\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10438\,
            I => \inst_midgetv_core.ADR_O_4\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__10435\,
            I => \inst_midgetv_core.ADR_O_4\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__10426\,
            I => \N__10423\
        );

    \I__2261\ : CascadeBuf
    port map (
            O => \N__10423\,
            I => \N__10420\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__10420\,
            I => \N__10417\
        );

    \I__2259\ : CascadeBuf
    port map (
            O => \N__10417\,
            I => \N__10414\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__10414\,
            I => \N__10411\
        );

    \I__2257\ : CascadeBuf
    port map (
            O => \N__10411\,
            I => \N__10408\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__10408\,
            I => \N__10405\
        );

    \I__2255\ : CascadeBuf
    port map (
            O => \N__10405\,
            I => \N__10402\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__10402\,
            I => \N__10399\
        );

    \I__2253\ : CascadeBuf
    port map (
            O => \N__10399\,
            I => \N__10396\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__10396\,
            I => \N__10393\
        );

    \I__2251\ : CascadeBuf
    port map (
            O => \N__10393\,
            I => \N__10390\
        );

    \I__2250\ : CascadeMux
    port map (
            O => \N__10390\,
            I => \N__10387\
        );

    \I__2249\ : CascadeBuf
    port map (
            O => \N__10387\,
            I => \N__10384\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__10384\,
            I => \N__10381\
        );

    \I__2247\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10378\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__10378\,
            I => \N__10375\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__10375\,
            I => \N__10372\
        );

    \I__2244\ : Span4Mux_v
    port map (
            O => \N__10372\,
            I => \N__10369\
        );

    \I__2243\ : Span4Mux_v
    port map (
            O => \N__10369\,
            I => \N__10366\
        );

    \I__2242\ : Span4Mux_v
    port map (
            O => \N__10366\,
            I => \N__10363\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__10363\,
            I => \inst_midgetv_core.Wai_2\
        );

    \I__2240\ : InMux
    port map (
            O => \N__10360\,
            I => \N__10357\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__10357\,
            I => \N__10351\
        );

    \I__2238\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10348\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10355\,
            I => \N__10345\
        );

    \I__2236\ : InMux
    port map (
            O => \N__10354\,
            I => \N__10342\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__10351\,
            I => \inst_midgetv_core.ADR_O_5\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__10348\,
            I => \inst_midgetv_core.ADR_O_5\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__10345\,
            I => \inst_midgetv_core.ADR_O_5\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__10342\,
            I => \inst_midgetv_core.ADR_O_5\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__10333\,
            I => \N__10330\
        );

    \I__2230\ : CascadeBuf
    port map (
            O => \N__10330\,
            I => \N__10327\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__10327\,
            I => \N__10324\
        );

    \I__2228\ : CascadeBuf
    port map (
            O => \N__10324\,
            I => \N__10321\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__10321\,
            I => \N__10318\
        );

    \I__2226\ : CascadeBuf
    port map (
            O => \N__10318\,
            I => \N__10315\
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__10315\,
            I => \N__10312\
        );

    \I__2224\ : CascadeBuf
    port map (
            O => \N__10312\,
            I => \N__10309\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__10309\,
            I => \N__10306\
        );

    \I__2222\ : CascadeBuf
    port map (
            O => \N__10306\,
            I => \N__10303\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__10303\,
            I => \N__10300\
        );

    \I__2220\ : CascadeBuf
    port map (
            O => \N__10300\,
            I => \N__10297\
        );

    \I__2219\ : CascadeMux
    port map (
            O => \N__10297\,
            I => \N__10294\
        );

    \I__2218\ : CascadeBuf
    port map (
            O => \N__10294\,
            I => \N__10291\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__10291\,
            I => \N__10288\
        );

    \I__2216\ : InMux
    port map (
            O => \N__10288\,
            I => \N__10285\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__10285\,
            I => \N__10282\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__10282\,
            I => \N__10279\
        );

    \I__2213\ : Sp12to4
    port map (
            O => \N__10279\,
            I => \N__10276\
        );

    \I__2212\ : Span12Mux_s8_h
    port map (
            O => \N__10276\,
            I => \N__10273\
        );

    \I__2211\ : Odrv12
    port map (
            O => \N__10273\,
            I => \inst_midgetv_core.Wai_3\
        );

    \I__2210\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10266\
        );

    \I__2209\ : InMux
    port map (
            O => \N__10269\,
            I => \N__10263\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__10266\,
            I => \N__10259\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__10263\,
            I => \N__10256\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__10262\,
            I => \N__10253\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__10259\,
            I => \N__10248\
        );

    \I__2204\ : Span4Mux_v
    port map (
            O => \N__10256\,
            I => \N__10248\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10245\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__10248\,
            I => \inst_midgetv_core.INSTR_11\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__10245\,
            I => \inst_midgetv_core.INSTR_11\
        );

    \I__2200\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10237\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__10237\,
            I => \N__10234\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__10234\,
            I => \N__10231\
        );

    \I__2197\ : Span4Mux_h
    port map (
            O => \N__10231\,
            I => \N__10225\
        );

    \I__2196\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10222\
        );

    \I__2195\ : InMux
    port map (
            O => \N__10229\,
            I => \N__10217\
        );

    \I__2194\ : InMux
    port map (
            O => \N__10228\,
            I => \N__10217\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__10225\,
            I => \inst_midgetv_core.ADR_O_6\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__10222\,
            I => \inst_midgetv_core.ADR_O_6\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__10217\,
            I => \inst_midgetv_core.ADR_O_6\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__10210\,
            I => \N__10207\
        );

    \I__2189\ : CascadeBuf
    port map (
            O => \N__10207\,
            I => \N__10204\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__10204\,
            I => \N__10201\
        );

    \I__2187\ : CascadeBuf
    port map (
            O => \N__10201\,
            I => \N__10198\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__10198\,
            I => \N__10195\
        );

    \I__2185\ : CascadeBuf
    port map (
            O => \N__10195\,
            I => \N__10192\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__10192\,
            I => \N__10189\
        );

    \I__2183\ : CascadeBuf
    port map (
            O => \N__10189\,
            I => \N__10186\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__10186\,
            I => \N__10183\
        );

    \I__2181\ : CascadeBuf
    port map (
            O => \N__10183\,
            I => \N__10180\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__10180\,
            I => \N__10177\
        );

    \I__2179\ : CascadeBuf
    port map (
            O => \N__10177\,
            I => \N__10174\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__10174\,
            I => \N__10171\
        );

    \I__2177\ : CascadeBuf
    port map (
            O => \N__10171\,
            I => \N__10168\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__10168\,
            I => \N__10165\
        );

    \I__2175\ : InMux
    port map (
            O => \N__10165\,
            I => \N__10162\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__10162\,
            I => \N__10159\
        );

    \I__2173\ : Span4Mux_s3_v
    port map (
            O => \N__10159\,
            I => \N__10156\
        );

    \I__2172\ : Sp12to4
    port map (
            O => \N__10156\,
            I => \N__10153\
        );

    \I__2171\ : Span12Mux_s8_h
    port map (
            O => \N__10153\,
            I => \N__10150\
        );

    \I__2170\ : Span12Mux_v
    port map (
            O => \N__10150\,
            I => \N__10147\
        );

    \I__2169\ : Odrv12
    port map (
            O => \N__10147\,
            I => \inst_midgetv_core.Wai_4\
        );

    \I__2168\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10139\
        );

    \I__2167\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10136\
        );

    \I__2166\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10133\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__10139\,
            I => \N__10129\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__10136\,
            I => \N__10126\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__10133\,
            I => \N__10123\
        );

    \I__2162\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10120\
        );

    \I__2161\ : Odrv12
    port map (
            O => \N__10129\,
            I => \inst_midgetv_core.ADR_O_7\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__10126\,
            I => \inst_midgetv_core.ADR_O_7\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__10123\,
            I => \inst_midgetv_core.ADR_O_7\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__10120\,
            I => \inst_midgetv_core.ADR_O_7\
        );

    \I__2157\ : InMux
    port map (
            O => \N__10111\,
            I => \inst_midgetv_core.inst_wai.genblk1_waicy4\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__10108\,
            I => \N__10105\
        );

    \I__2155\ : CascadeBuf
    port map (
            O => \N__10105\,
            I => \N__10102\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__10102\,
            I => \N__10099\
        );

    \I__2153\ : CascadeBuf
    port map (
            O => \N__10099\,
            I => \N__10096\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__10096\,
            I => \N__10093\
        );

    \I__2151\ : CascadeBuf
    port map (
            O => \N__10093\,
            I => \N__10090\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__10090\,
            I => \N__10087\
        );

    \I__2149\ : CascadeBuf
    port map (
            O => \N__10087\,
            I => \N__10084\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__10084\,
            I => \N__10081\
        );

    \I__2147\ : CascadeBuf
    port map (
            O => \N__10081\,
            I => \N__10078\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__10078\,
            I => \N__10075\
        );

    \I__2145\ : CascadeBuf
    port map (
            O => \N__10075\,
            I => \N__10072\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__10072\,
            I => \N__10069\
        );

    \I__2143\ : CascadeBuf
    port map (
            O => \N__10069\,
            I => \N__10066\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__10066\,
            I => \N__10063\
        );

    \I__2141\ : InMux
    port map (
            O => \N__10063\,
            I => \N__10060\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__10060\,
            I => \N__10057\
        );

    \I__2139\ : Span4Mux_s2_v
    port map (
            O => \N__10057\,
            I => \N__10054\
        );

    \I__2138\ : Sp12to4
    port map (
            O => \N__10054\,
            I => \N__10051\
        );

    \I__2137\ : Span12Mux_v
    port map (
            O => \N__10051\,
            I => \N__10048\
        );

    \I__2136\ : Odrv12
    port map (
            O => \N__10048\,
            I => \inst_midgetv_core.Wai_5\
        );

    \I__2135\ : InMux
    port map (
            O => \N__10045\,
            I => \N__10042\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__10042\,
            I => \inst_midgetv_core.inst_wai.genblk1_preWai0\
        );

    \I__2133\ : InMux
    port map (
            O => \N__10039\,
            I => \N__10034\
        );

    \I__2132\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10031\
        );

    \I__2131\ : InMux
    port map (
            O => \N__10037\,
            I => \N__10028\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__10034\,
            I => \N__10025\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__10031\,
            I => \N__10020\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__10028\,
            I => \N__10020\
        );

    \I__2127\ : Span4Mux_v
    port map (
            O => \N__10025\,
            I => \N__10014\
        );

    \I__2126\ : Span4Mux_v
    port map (
            O => \N__10020\,
            I => \N__10014\
        );

    \I__2125\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10011\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__10014\,
            I => \inst_midgetv_core.INSTR_7\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__10011\,
            I => \inst_midgetv_core.INSTR_7\
        );

    \I__2122\ : InMux
    port map (
            O => \N__10006\,
            I => \N__10003\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__10003\,
            I => \N__10000\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__10000\,
            I => \N__9997\
        );

    \I__2119\ : Span4Mux_h
    port map (
            O => \N__9997\,
            I => \N__9994\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__9994\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm0a\
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__9991\,
            I => \N__9988\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9984\
        );

    \I__2115\ : InMux
    port map (
            O => \N__9987\,
            I => \N__9981\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9984\,
            I => \N__9977\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__9981\,
            I => \N__9974\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9971\
        );

    \I__2111\ : Span4Mux_h
    port map (
            O => \N__9977\,
            I => \N__9968\
        );

    \I__2110\ : Span4Mux_h
    port map (
            O => \N__9974\,
            I => \N__9965\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__9971\,
            I => \N__9962\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__9968\,
            I => \inst_midgetv_core.INSTR_9\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__9965\,
            I => \inst_midgetv_core.INSTR_9\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__9962\,
            I => \inst_midgetv_core.INSTR_9\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9955\,
            I => \N__9952\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9952\,
            I => \N__9949\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__9949\,
            I => \N__9946\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__9946\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm2a\
        );

    \I__2101\ : CEMux
    port map (
            O => \N__9943\,
            I => \N__9939\
        );

    \I__2100\ : CEMux
    port map (
            O => \N__9942\,
            I => \N__9936\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9939\,
            I => \N__9933\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__9936\,
            I => \N__9930\
        );

    \I__2097\ : Span4Mux_v
    port map (
            O => \N__9933\,
            I => \N__9927\
        );

    \I__2096\ : Span4Mux_h
    port map (
            O => \N__9930\,
            I => \N__9924\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__9927\,
            I => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.we\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__9924\,
            I => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.we\
        );

    \I__2093\ : CEMux
    port map (
            O => \N__9919\,
            I => \N__9915\
        );

    \I__2092\ : CEMux
    port map (
            O => \N__9918\,
            I => \N__9912\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__9915\,
            I => \N__9908\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9912\,
            I => \N__9905\
        );

    \I__2089\ : CEMux
    port map (
            O => \N__9911\,
            I => \N__9902\
        );

    \I__2088\ : Span4Mux_v
    port map (
            O => \N__9908\,
            I => \N__9895\
        );

    \I__2087\ : Span4Mux_v
    port map (
            O => \N__9905\,
            I => \N__9892\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9902\,
            I => \N__9889\
        );

    \I__2085\ : CEMux
    port map (
            O => \N__9901\,
            I => \N__9886\
        );

    \I__2084\ : CEMux
    port map (
            O => \N__9900\,
            I => \N__9883\
        );

    \I__2083\ : CEMux
    port map (
            O => \N__9899\,
            I => \N__9880\
        );

    \I__2082\ : CEMux
    port map (
            O => \N__9898\,
            I => \N__9877\
        );

    \I__2081\ : Span4Mux_h
    port map (
            O => \N__9895\,
            I => \N__9873\
        );

    \I__2080\ : Span4Mux_h
    port map (
            O => \N__9892\,
            I => \N__9868\
        );

    \I__2079\ : Span4Mux_h
    port map (
            O => \N__9889\,
            I => \N__9868\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9886\,
            I => \N__9865\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__9883\,
            I => \N__9862\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9880\,
            I => \N__9859\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__9877\,
            I => \N__9856\
        );

    \I__2074\ : CEMux
    port map (
            O => \N__9876\,
            I => \N__9853\
        );

    \I__2073\ : Sp12to4
    port map (
            O => \N__9873\,
            I => \N__9850\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__9868\,
            I => \N__9847\
        );

    \I__2071\ : Span4Mux_h
    port map (
            O => \N__9865\,
            I => \N__9844\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__9862\,
            I => \N__9841\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__9859\,
            I => \N__9838\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__9856\,
            I => \N__9833\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__9853\,
            I => \N__9833\
        );

    \I__2066\ : Span12Mux_v
    port map (
            O => \N__9850\,
            I => \N__9830\
        );

    \I__2065\ : Span4Mux_h
    port map (
            O => \N__9847\,
            I => \N__9827\
        );

    \I__2064\ : Span4Mux_h
    port map (
            O => \N__9844\,
            I => \N__9824\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__9841\,
            I => \N__9817\
        );

    \I__2062\ : Span4Mux_h
    port map (
            O => \N__9838\,
            I => \N__9817\
        );

    \I__2061\ : Span4Mux_v
    port map (
            O => \N__9833\,
            I => \N__9817\
        );

    \I__2060\ : Odrv12
    port map (
            O => \N__9830\,
            I => \inst_midgetv_core.is_valid_instrhigh\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__9827\,
            I => \inst_midgetv_core.is_valid_instrhigh\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__9824\,
            I => \inst_midgetv_core.is_valid_instrhigh\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__9817\,
            I => \inst_midgetv_core.is_valid_instrhigh\
        );

    \I__2056\ : CEMux
    port map (
            O => \N__9808\,
            I => \N__9803\
        );

    \I__2055\ : SRMux
    port map (
            O => \N__9807\,
            I => \N__9800\
        );

    \I__2054\ : SRMux
    port map (
            O => \N__9806\,
            I => \N__9797\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9803\,
            I => \N__9794\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9800\,
            I => \N__9791\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9797\,
            I => \N__9788\
        );

    \I__2050\ : Span4Mux_h
    port map (
            O => \N__9794\,
            I => \N__9785\
        );

    \I__2049\ : Span4Mux_v
    port map (
            O => \N__9791\,
            I => \N__9782\
        );

    \I__2048\ : Span4Mux_h
    port map (
            O => \N__9788\,
            I => \N__9779\
        );

    \I__2047\ : Odrv4
    port map (
            O => \N__9785\,
            I => \inst_midgetv_core.progress_ucode\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__9782\,
            I => \inst_midgetv_core.progress_ucode\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__9779\,
            I => \inst_midgetv_core.progress_ucode\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__9772\,
            I => \N__9769\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9766\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9766\,
            I => \N__9763\
        );

    \I__2041\ : Span4Mux_h
    port map (
            O => \N__9763\,
            I => \N__9760\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__9760\,
            I => \inst_midgetv_core.rinx_0\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9757\,
            I => \N__9754\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9754\,
            I => \N__9751\
        );

    \I__2037\ : Odrv12
    port map (
            O => \N__9751\,
            I => \inst_midgetv_core.inst_ucodepc.n5624\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9745\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9745\,
            I => \inst_midgetv_core.sa33\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9739\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9739\,
            I => \inst_midgetv_core.inst_progressctrl.n4\
        );

    \I__2032\ : CEMux
    port map (
            O => \N__9736\,
            I => \N__9732\
        );

    \I__2031\ : CEMux
    port map (
            O => \N__9735\,
            I => \N__9729\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9732\,
            I => \N__9721\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9729\,
            I => \N__9721\
        );

    \I__2028\ : CEMux
    port map (
            O => \N__9728\,
            I => \N__9718\
        );

    \I__2027\ : CEMux
    port map (
            O => \N__9727\,
            I => \N__9715\
        );

    \I__2026\ : CEMux
    port map (
            O => \N__9726\,
            I => \N__9712\
        );

    \I__2025\ : Span4Mux_v
    port map (
            O => \N__9721\,
            I => \N__9707\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9718\,
            I => \N__9707\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9715\,
            I => \N__9704\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__9712\,
            I => \N__9701\
        );

    \I__2021\ : Span4Mux_v
    port map (
            O => \N__9707\,
            I => \N__9698\
        );

    \I__2020\ : Span4Mux_h
    port map (
            O => \N__9704\,
            I => \N__9695\
        );

    \I__2019\ : Span4Mux_v
    port map (
            O => \N__9701\,
            I => \N__9690\
        );

    \I__2018\ : Span4Mux_h
    port map (
            O => \N__9698\,
            I => \N__9690\
        );

    \I__2017\ : Span4Mux_h
    port map (
            O => \N__9695\,
            I => \N__9687\
        );

    \I__2016\ : Span4Mux_h
    port map (
            O => \N__9690\,
            I => \N__9684\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__9687\,
            I => \inst_midgetv_core.enaQ\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__9684\,
            I => \inst_midgetv_core.enaQ\
        );

    \I__2013\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9676\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__9676\,
            I => \N__9673\
        );

    \I__2011\ : Span4Mux_h
    port map (
            O => \N__9673\,
            I => \N__9670\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__9670\,
            I => \inst_midgetv_core.sa00\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__9667\,
            I => \N__9664\
        );

    \I__2008\ : CascadeBuf
    port map (
            O => \N__9664\,
            I => \N__9661\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__9661\,
            I => \N__9658\
        );

    \I__2006\ : CascadeBuf
    port map (
            O => \N__9658\,
            I => \N__9655\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__9655\,
            I => \N__9652\
        );

    \I__2004\ : CascadeBuf
    port map (
            O => \N__9652\,
            I => \N__9649\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__9649\,
            I => \N__9646\
        );

    \I__2002\ : CascadeBuf
    port map (
            O => \N__9646\,
            I => \N__9643\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__9643\,
            I => \N__9640\
        );

    \I__2000\ : CascadeBuf
    port map (
            O => \N__9640\,
            I => \N__9637\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__9637\,
            I => \N__9634\
        );

    \I__1998\ : CascadeBuf
    port map (
            O => \N__9634\,
            I => \N__9631\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__9631\,
            I => \N__9628\
        );

    \I__1996\ : CascadeBuf
    port map (
            O => \N__9628\,
            I => \N__9625\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__9625\,
            I => \N__9622\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9622\,
            I => \N__9619\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9619\,
            I => \N__9616\
        );

    \I__1992\ : Span4Mux_s3_v
    port map (
            O => \N__9616\,
            I => \N__9613\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__9613\,
            I => \N__9610\
        );

    \I__1990\ : Span4Mux_v
    port map (
            O => \N__9610\,
            I => \N__9607\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__9607\,
            I => \N__9604\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__9604\,
            I => \inst_midgetv_core.Wai_0\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__9601\,
            I => \N__9596\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9591\
        );

    \I__1985\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9591\
        );

    \I__1984\ : InMux
    port map (
            O => \N__9596\,
            I => \N__9588\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__9591\,
            I => \N__9585\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__9588\,
            I => \N__9582\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__9585\,
            I => \N__9579\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__9582\,
            I => \inst_midgetv_core.ADR_O_14\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__9579\,
            I => \inst_midgetv_core.ADR_O_14\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__9574\,
            I => \inst_midgetv_core.Di_14_cascade_\
        );

    \I__1977\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9568\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__9568\,
            I => \N__9565\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__9565\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_14\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__9562\,
            I => \N__9559\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9559\,
            I => \N__9556\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__9556\,
            I => \N__9553\
        );

    \I__1971\ : Span4Mux_v
    port map (
            O => \N__9553\,
            I => \N__9550\
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__9550\,
            I => \inst_midgetv_core.DAT_O_15\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__9547\,
            I => \N__9544\
        );

    \I__1968\ : InMux
    port map (
            O => \N__9544\,
            I => \N__9539\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9534\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9542\,
            I => \N__9534\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9539\,
            I => \N__9531\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__9534\,
            I => \N__9528\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__9531\,
            I => \N__9523\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__9528\,
            I => \N__9523\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__9523\,
            I => \inst_midgetv_core.ADR_O_15\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__9520\,
            I => \inst_midgetv_core.Di_15_cascade_\
        );

    \I__1959\ : InMux
    port map (
            O => \N__9517\,
            I => \N__9514\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__9514\,
            I => \N__9511\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__9511\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_15\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__9508\,
            I => \N__9503\
        );

    \I__1955\ : InMux
    port map (
            O => \N__9507\,
            I => \N__9500\
        );

    \I__1954\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9497\
        );

    \I__1953\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9494\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__9500\,
            I => \N__9489\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__9497\,
            I => \N__9489\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__9494\,
            I => \N__9484\
        );

    \I__1949\ : Span4Mux_h
    port map (
            O => \N__9489\,
            I => \N__9484\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__9484\,
            I => \inst_midgetv_core.ADR_O_17\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__9481\,
            I => \N__9478\
        );

    \I__1946\ : InMux
    port map (
            O => \N__9478\,
            I => \N__9475\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__9475\,
            I => \N__9472\
        );

    \I__1944\ : Span4Mux_h
    port map (
            O => \N__9472\,
            I => \N__9469\
        );

    \I__1943\ : Span4Mux_v
    port map (
            O => \N__9469\,
            I => \N__9466\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__9466\,
            I => \inst_midgetv_core.DAT_O_16\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9463\,
            I => \N__9446\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9462\,
            I => \N__9446\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9446\
        );

    \I__1938\ : InMux
    port map (
            O => \N__9460\,
            I => \N__9446\
        );

    \I__1937\ : InMux
    port map (
            O => \N__9459\,
            I => \N__9436\
        );

    \I__1936\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9436\
        );

    \I__1935\ : InMux
    port map (
            O => \N__9457\,
            I => \N__9436\
        );

    \I__1934\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9436\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__9455\,
            I => \N__9432\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__9446\,
            I => \N__9415\
        );

    \I__1931\ : InMux
    port map (
            O => \N__9445\,
            I => \N__9412\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__9436\,
            I => \N__9409\
        );

    \I__1929\ : InMux
    port map (
            O => \N__9435\,
            I => \N__9400\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9432\,
            I => \N__9400\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9400\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9400\
        );

    \I__1925\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9391\
        );

    \I__1924\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9391\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9391\
        );

    \I__1922\ : InMux
    port map (
            O => \N__9426\,
            I => \N__9391\
        );

    \I__1921\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9382\
        );

    \I__1920\ : InMux
    port map (
            O => \N__9424\,
            I => \N__9382\
        );

    \I__1919\ : InMux
    port map (
            O => \N__9423\,
            I => \N__9382\
        );

    \I__1918\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9382\
        );

    \I__1917\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9366\
        );

    \I__1916\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9366\
        );

    \I__1915\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9366\
        );

    \I__1914\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9366\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__9415\,
            I => \N__9361\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__9412\,
            I => \N__9361\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__9409\,
            I => \N__9352\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__9400\,
            I => \N__9352\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__9391\,
            I => \N__9352\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__9382\,
            I => \N__9352\
        );

    \I__1907\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9345\
        );

    \I__1906\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9345\
        );

    \I__1905\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9345\
        );

    \I__1904\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9336\
        );

    \I__1903\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9336\
        );

    \I__1902\ : InMux
    port map (
            O => \N__9376\,
            I => \N__9336\
        );

    \I__1901\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9336\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__9366\,
            I => \inst_midgetv_core.inst_mimux.genblk1_sa00mod\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__9361\,
            I => \inst_midgetv_core.inst_mimux.genblk1_sa00mod\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__9352\,
            I => \inst_midgetv_core.inst_mimux.genblk1_sa00mod\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__9345\,
            I => \inst_midgetv_core.inst_mimux.genblk1_sa00mod\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__9336\,
            I => \inst_midgetv_core.inst_mimux.genblk1_sa00mod\
        );

    \I__1895\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9318\
        );

    \I__1894\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9318\
        );

    \I__1893\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9315\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__9318\,
            I => \N__9312\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__9315\,
            I => \N__9307\
        );

    \I__1890\ : Span4Mux_h
    port map (
            O => \N__9312\,
            I => \N__9307\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__9307\,
            I => \inst_midgetv_core.ADR_O_16\
        );

    \I__1888\ : InMux
    port map (
            O => \N__9304\,
            I => \N__9284\
        );

    \I__1887\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9284\
        );

    \I__1886\ : InMux
    port map (
            O => \N__9302\,
            I => \N__9284\
        );

    \I__1885\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9284\
        );

    \I__1884\ : InMux
    port map (
            O => \N__9300\,
            I => \N__9275\
        );

    \I__1883\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9275\
        );

    \I__1882\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9275\
        );

    \I__1881\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9275\
        );

    \I__1880\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9268\
        );

    \I__1879\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9268\
        );

    \I__1878\ : InMux
    port map (
            O => \N__9294\,
            I => \N__9268\
        );

    \I__1877\ : InMux
    port map (
            O => \N__9293\,
            I => \N__9265\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__9284\,
            I => \N__9244\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__9275\,
            I => \N__9237\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__9268\,
            I => \N__9237\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__9265\,
            I => \N__9237\
        );

    \I__1872\ : InMux
    port map (
            O => \N__9264\,
            I => \N__9230\
        );

    \I__1871\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9230\
        );

    \I__1870\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9230\
        );

    \I__1869\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9221\
        );

    \I__1868\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9221\
        );

    \I__1867\ : InMux
    port map (
            O => \N__9259\,
            I => \N__9221\
        );

    \I__1866\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9221\
        );

    \I__1865\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9212\
        );

    \I__1864\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9212\
        );

    \I__1863\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9212\
        );

    \I__1862\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9212\
        );

    \I__1861\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9209\
        );

    \I__1860\ : InMux
    port map (
            O => \N__9252\,
            I => \N__9202\
        );

    \I__1859\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9202\
        );

    \I__1858\ : InMux
    port map (
            O => \N__9250\,
            I => \N__9202\
        );

    \I__1857\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9199\
        );

    \I__1856\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9192\
        );

    \I__1855\ : InMux
    port map (
            O => \N__9247\,
            I => \N__9192\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__9244\,
            I => \N__9189\
        );

    \I__1853\ : Span4Mux_v
    port map (
            O => \N__9237\,
            I => \N__9180\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__9230\,
            I => \N__9180\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__9221\,
            I => \N__9180\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__9212\,
            I => \N__9180\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__9209\,
            I => \N__9173\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__9202\,
            I => \N__9173\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__9199\,
            I => \N__9173\
        );

    \I__1846\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9168\
        );

    \I__1845\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9168\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__9192\,
            I => \N__9165\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__9189\,
            I => \N__9162\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__9180\,
            I => \N__9159\
        );

    \I__1841\ : Span4Mux_v
    port map (
            O => \N__9173\,
            I => \N__9154\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__9168\,
            I => \N__9154\
        );

    \I__1839\ : Span4Mux_h
    port map (
            O => \N__9165\,
            I => \N__9151\
        );

    \I__1838\ : Span4Mux_h
    port map (
            O => \N__9162\,
            I => \N__9148\
        );

    \I__1837\ : Span4Mux_h
    port map (
            O => \N__9159\,
            I => \N__9145\
        );

    \I__1836\ : Span4Mux_v
    port map (
            O => \N__9154\,
            I => \N__9142\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__9151\,
            I => \N__9139\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__9148\,
            I => \inst_midgetv_core.s_alu_1\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__9145\,
            I => \inst_midgetv_core.s_alu_1\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__9142\,
            I => \inst_midgetv_core.s_alu_1\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__9139\,
            I => \inst_midgetv_core.s_alu_1\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__9130\,
            I => \inst_midgetv_core.Di_16_cascade_\
        );

    \I__1829\ : InMux
    port map (
            O => \N__9127\,
            I => \N__9100\
        );

    \I__1828\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9100\
        );

    \I__1827\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9100\
        );

    \I__1826\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9100\
        );

    \I__1825\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9093\
        );

    \I__1824\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9093\
        );

    \I__1823\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9093\
        );

    \I__1822\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9090\
        );

    \I__1821\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9076\
        );

    \I__1820\ : InMux
    port map (
            O => \N__9118\,
            I => \N__9076\
        );

    \I__1819\ : InMux
    port map (
            O => \N__9117\,
            I => \N__9067\
        );

    \I__1818\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9067\
        );

    \I__1817\ : InMux
    port map (
            O => \N__9115\,
            I => \N__9067\
        );

    \I__1816\ : InMux
    port map (
            O => \N__9114\,
            I => \N__9067\
        );

    \I__1815\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9058\
        );

    \I__1814\ : InMux
    port map (
            O => \N__9112\,
            I => \N__9058\
        );

    \I__1813\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9058\
        );

    \I__1812\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9058\
        );

    \I__1811\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9055\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__9100\,
            I => \N__9052\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__9093\,
            I => \N__9049\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__9090\,
            I => \N__9046\
        );

    \I__1807\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9037\
        );

    \I__1806\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9037\
        );

    \I__1805\ : InMux
    port map (
            O => \N__9087\,
            I => \N__9037\
        );

    \I__1804\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9037\
        );

    \I__1803\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9032\
        );

    \I__1802\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9032\
        );

    \I__1801\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9025\
        );

    \I__1800\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9025\
        );

    \I__1799\ : InMux
    port map (
            O => \N__9081\,
            I => \N__9025\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__9076\,
            I => \N__9016\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__9067\,
            I => \N__9016\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__9058\,
            I => \N__9016\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__9055\,
            I => \N__9016\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__9052\,
            I => \N__9009\
        );

    \I__1793\ : Span4Mux_v
    port map (
            O => \N__9049\,
            I => \N__8998\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__9046\,
            I => \N__8998\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__9037\,
            I => \N__8998\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__9032\,
            I => \N__8998\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__9025\,
            I => \N__8998\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__9016\,
            I => \N__8995\
        );

    \I__1787\ : InMux
    port map (
            O => \N__9015\,
            I => \N__8986\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9014\,
            I => \N__8986\
        );

    \I__1785\ : InMux
    port map (
            O => \N__9013\,
            I => \N__8986\
        );

    \I__1784\ : InMux
    port map (
            O => \N__9012\,
            I => \N__8986\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__9009\,
            I => \N__8983\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__8998\,
            I => \N__8980\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__8995\,
            I => \N__8975\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8986\,
            I => \N__8975\
        );

    \I__1779\ : Span4Mux_h
    port map (
            O => \N__8983\,
            I => \N__8972\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__8980\,
            I => \N__8967\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__8975\,
            I => \N__8967\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__8972\,
            I => \inst_midgetv_core.s_alu_0\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__8967\,
            I => \inst_midgetv_core.s_alu_0\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__8962\,
            I => \N__8959\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8956\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8956\,
            I => \N__8953\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__8953\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_16\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8947\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8947\,
            I => \N__8944\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__8944\,
            I => \N__8940\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8943\,
            I => \N__8936\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__8940\,
            I => \N__8932\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8929\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8936\,
            I => \N__8926\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8923\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__8932\,
            I => \N__8918\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8929\,
            I => \N__8918\
        );

    \I__1760\ : Span4Mux_h
    port map (
            O => \N__8926\,
            I => \N__8915\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8923\,
            I => \inst_midgetv_core.B_30\
        );

    \I__1758\ : Odrv4
    port map (
            O => \N__8918\,
            I => \inst_midgetv_core.B_30\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__8915\,
            I => \inst_midgetv_core.B_30\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8905\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__8905\,
            I => \N__8902\
        );

    \I__1754\ : Odrv12
    port map (
            O => \N__8902\,
            I => \inst_midgetv_core.sa29\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8896\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8896\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk1_illegal_rs1_rd_N_300\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8890\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8890\,
            I => \uart_ACK_O\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__8887\,
            I => \N__8883\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8880\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8877\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8880\,
            I => \rDee_8\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8877\,
            I => \rDee_8\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__8872\,
            I => \N__8869\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8863\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8858\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8858\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8855\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8863\,
            I => \N__8850\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8858\,
            I => \N__8850\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__8855\,
            I => \N__8846\
        );

    \I__1736\ : Span4Mux_h
    port map (
            O => \N__8850\,
            I => \N__8843\
        );

    \I__1735\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8840\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__8846\,
            I => \inst_midgetv_core.FUNC7_6\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__8843\,
            I => \inst_midgetv_core.FUNC7_6\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8840\,
            I => \inst_midgetv_core.FUNC7_6\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8830\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__8830\,
            I => \N__8826\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8829\,
            I => \N__8822\
        );

    \I__1728\ : Span4Mux_h
    port map (
            O => \N__8826\,
            I => \N__8819\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8816\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__8822\,
            I => \N__8813\
        );

    \I__1725\ : Span4Mux_h
    port map (
            O => \N__8819\,
            I => \N__8808\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8816\,
            I => \N__8808\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__8813\,
            I => \N__8805\
        );

    \I__1722\ : Span4Mux_v
    port map (
            O => \N__8808\,
            I => \N__8802\
        );

    \I__1721\ : Odrv4
    port map (
            O => \N__8805\,
            I => \inst_midgetv_core.FUNC7_1\
        );

    \I__1720\ : Odrv4
    port map (
            O => \N__8802\,
            I => \inst_midgetv_core.FUNC7_1\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8797\,
            I => \N__8792\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8796\,
            I => \N__8789\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__8795\,
            I => \N__8786\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8792\,
            I => \N__8783\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8789\,
            I => \N__8780\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8777\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__8783\,
            I => \N__8772\
        );

    \I__1712\ : Span4Mux_v
    port map (
            O => \N__8780\,
            I => \N__8772\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8777\,
            I => \N__8769\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__8772\,
            I => \inst_midgetv_core.FUNC7_3\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__8769\,
            I => \inst_midgetv_core.FUNC7_3\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8761\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__8761\,
            I => \N__8757\
        );

    \I__1706\ : InMux
    port map (
            O => \N__8760\,
            I => \N__8753\
        );

    \I__1705\ : Span4Mux_v
    port map (
            O => \N__8757\,
            I => \N__8750\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8746\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__8753\,
            I => \N__8743\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__8750\,
            I => \N__8740\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8749\,
            I => \N__8737\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8746\,
            I => \N__8734\
        );

    \I__1699\ : Span4Mux_h
    port map (
            O => \N__8743\,
            I => \N__8731\
        );

    \I__1698\ : Sp12to4
    port map (
            O => \N__8740\,
            I => \N__8728\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8737\,
            I => \N__8723\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__8734\,
            I => \N__8723\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__8731\,
            I => \inst_midgetv_core.FUNC7_0\
        );

    \I__1694\ : Odrv12
    port map (
            O => \N__8728\,
            I => \inst_midgetv_core.FUNC7_0\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__8723\,
            I => \inst_midgetv_core.FUNC7_0\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8716\,
            I => \N__8713\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__8713\,
            I => \N__8710\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__8710\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n12\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8704\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8704\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n17\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__8701\,
            I => \N__8698\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8695\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8695\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n16\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__8692\,
            I => \N__8689\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8686\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__8686\,
            I => \N__8683\
        );

    \I__1681\ : Span4Mux_h
    port map (
            O => \N__8683\,
            I => \N__8680\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__8680\,
            I => \inst_midgetv_core.DAT_O_13\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8672\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8667\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8667\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__8672\,
            I => \N__8660\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8667\,
            I => \N__8657\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8654\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8665\,
            I => \N__8651\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8646\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8646\
        );

    \I__1670\ : Span4Mux_h
    port map (
            O => \N__8660\,
            I => \N__8643\
        );

    \I__1669\ : Span4Mux_h
    port map (
            O => \N__8657\,
            I => \N__8640\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__8654\,
            I => \N__8637\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8651\,
            I => \N__8632\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8646\,
            I => \N__8632\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__8643\,
            I => \inst_midgetv_core.INSTR_13\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__8640\,
            I => \inst_midgetv_core.INSTR_13\
        );

    \I__1663\ : Odrv12
    port map (
            O => \N__8637\,
            I => \inst_midgetv_core.INSTR_13\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__8632\,
            I => \inst_midgetv_core.INSTR_13\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__8623\,
            I => \inst_midgetv_core.Di_13_cascade_\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__8620\,
            I => \N__8616\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8613\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8610\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__8613\,
            I => \N__8607\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__8610\,
            I => \N__8601\
        );

    \I__1655\ : Span4Mux_h
    port map (
            O => \N__8607\,
            I => \N__8601\
        );

    \I__1654\ : InMux
    port map (
            O => \N__8606\,
            I => \N__8598\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__8601\,
            I => \inst_midgetv_core.ADR_O_13\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__8598\,
            I => \inst_midgetv_core.ADR_O_13\
        );

    \I__1651\ : InMux
    port map (
            O => \N__8593\,
            I => \N__8590\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8590\,
            I => \N__8587\
        );

    \I__1649\ : Odrv12
    port map (
            O => \N__8587\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_13\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__8584\,
            I => \N__8581\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8578\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__8578\,
            I => \N__8575\
        );

    \I__1645\ : Span4Mux_h
    port map (
            O => \N__8575\,
            I => \N__8572\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__8572\,
            I => \inst_midgetv_core.DAT_O_14\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8565\
        );

    \I__1642\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8562\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8565\,
            I => \N__8556\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__8562\,
            I => \N__8553\
        );

    \I__1639\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8550\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8560\,
            I => \N__8547\
        );

    \I__1637\ : InMux
    port map (
            O => \N__8559\,
            I => \N__8544\
        );

    \I__1636\ : Span4Mux_h
    port map (
            O => \N__8556\,
            I => \N__8541\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__8553\,
            I => \N__8538\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__8550\,
            I => \N__8535\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__8547\,
            I => \N__8530\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__8544\,
            I => \N__8530\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__8541\,
            I => \inst_midgetv_core.INSTR_14\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__8538\,
            I => \inst_midgetv_core.INSTR_14\
        );

    \I__1629\ : Odrv12
    port map (
            O => \N__8535\,
            I => \inst_midgetv_core.INSTR_14\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__8530\,
            I => \inst_midgetv_core.INSTR_14\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8518\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__8518\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n5605\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__8515\,
            I => \N__8507\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__8514\,
            I => \N__8504\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__8513\,
            I => \N__8501\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__8512\,
            I => \N__8498\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8493\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8510\,
            I => \N__8493\
        );

    \I__1619\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8490\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8485\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8485\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8498\,
            I => \N__8482\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__8493\,
            I => \inst_midgetv_core.INSTR_3\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__8490\,
            I => \inst_midgetv_core.INSTR_3\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__8485\,
            I => \inst_midgetv_core.INSTR_3\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8482\,
            I => \inst_midgetv_core.INSTR_3\
        );

    \I__1611\ : InMux
    port map (
            O => \N__8473\,
            I => \N__8470\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8470\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n8\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8462\
        );

    \I__1608\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8459\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8456\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__8462\,
            I => \N__8453\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__8459\,
            I => \N__8450\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__8456\,
            I => \N__8443\
        );

    \I__1603\ : Span4Mux_v
    port map (
            O => \N__8453\,
            I => \N__8443\
        );

    \I__1602\ : Span4Mux_h
    port map (
            O => \N__8450\,
            I => \N__8443\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__8443\,
            I => \inst_midgetv_core.FUNC7_2\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8440\,
            I => \N__8435\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8439\,
            I => \N__8432\
        );

    \I__1598\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8429\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__8435\,
            I => \N__8426\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__8432\,
            I => \N__8423\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8429\,
            I => \inst_midgetv_core.FUNC7_4\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__8426\,
            I => \inst_midgetv_core.FUNC7_4\
        );

    \I__1593\ : Odrv4
    port map (
            O => \N__8423\,
            I => \inst_midgetv_core.FUNC7_4\
        );

    \I__1592\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8411\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__8415\,
            I => \N__8408\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__8414\,
            I => \N__8405\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__8411\,
            I => \N__8401\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8397\
        );

    \I__1587\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8394\
        );

    \I__1586\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8391\
        );

    \I__1585\ : Span4Mux_v
    port map (
            O => \N__8401\,
            I => \N__8388\
        );

    \I__1584\ : InMux
    port map (
            O => \N__8400\,
            I => \N__8385\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__8397\,
            I => \N__8382\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__8394\,
            I => \N__8379\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__8391\,
            I => \N__8376\
        );

    \I__1580\ : Span4Mux_h
    port map (
            O => \N__8388\,
            I => \N__8371\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__8385\,
            I => \N__8371\
        );

    \I__1578\ : Span4Mux_h
    port map (
            O => \N__8382\,
            I => \N__8368\
        );

    \I__1577\ : Span12Mux_s10_h
    port map (
            O => \N__8379\,
            I => \N__8365\
        );

    \I__1576\ : Span4Mux_h
    port map (
            O => \N__8376\,
            I => \N__8362\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__8371\,
            I => \inst_midgetv_core.FUNC7_5\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__8368\,
            I => \inst_midgetv_core.FUNC7_5\
        );

    \I__1573\ : Odrv12
    port map (
            O => \N__8365\,
            I => \inst_midgetv_core.FUNC7_5\
        );

    \I__1572\ : Odrv4
    port map (
            O => \N__8362\,
            I => \inst_midgetv_core.FUNC7_5\
        );

    \I__1571\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8350\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__8350\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n497\
        );

    \I__1569\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8344\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__8344\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n11\
        );

    \I__1567\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8333\
        );

    \I__1566\ : InMux
    port map (
            O => \N__8340\,
            I => \N__8326\
        );

    \I__1565\ : InMux
    port map (
            O => \N__8339\,
            I => \N__8326\
        );

    \I__1564\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8326\
        );

    \I__1563\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8323\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__8336\,
            I => \N__8316\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__8333\,
            I => \N__8313\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8310\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__8323\,
            I => \N__8307\
        );

    \I__1558\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8302\
        );

    \I__1557\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8302\
        );

    \I__1556\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8297\
        );

    \I__1555\ : InMux
    port map (
            O => \N__8319\,
            I => \N__8297\
        );

    \I__1554\ : InMux
    port map (
            O => \N__8316\,
            I => \N__8294\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__8313\,
            I => \inst_midgetv_core.INSTR_5\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__8310\,
            I => \inst_midgetv_core.INSTR_5\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__8307\,
            I => \inst_midgetv_core.INSTR_5\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__8302\,
            I => \inst_midgetv_core.INSTR_5\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__8297\,
            I => \inst_midgetv_core.INSTR_5\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__8294\,
            I => \inst_midgetv_core.INSTR_5\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__8281\,
            I => \N__8278\
        );

    \I__1546\ : InMux
    port map (
            O => \N__8278\,
            I => \N__8274\
        );

    \I__1545\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8271\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__8274\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n2575\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__8271\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n2575\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__8266\,
            I => \N__8263\
        );

    \I__1541\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8260\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__8260\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk1_checkfunct7_N_281\
        );

    \I__1539\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8254\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__8254\,
            I => \N__8250\
        );

    \I__1537\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8247\
        );

    \I__1536\ : Span4Mux_h
    port map (
            O => \N__8250\,
            I => \N__8244\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__8247\,
            I => \N__8241\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__8244\,
            I => \inst_midgetv_core.raluF\
        );

    \I__1533\ : Odrv12
    port map (
            O => \N__8241\,
            I => \inst_midgetv_core.raluF\
        );

    \I__1532\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8233\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__8233\,
            I => \N__8230\
        );

    \I__1530\ : Span4Mux_h
    port map (
            O => \N__8230\,
            I => \N__8227\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__8227\,
            I => \inst_midgetv_core.is_brcond\
        );

    \I__1528\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8221\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__8221\,
            I => \N__8218\
        );

    \I__1526\ : Span4Mux_h
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__8215\,
            I => \inst_midgetv_core.rzcy32\
        );

    \I__1524\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8208\
        );

    \I__1523\ : InMux
    port map (
            O => \N__8211\,
            I => \N__8205\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__8208\,
            I => \N__8200\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__8205\,
            I => \N__8197\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__8204\,
            I => \N__8191\
        );

    \I__1519\ : InMux
    port map (
            O => \N__8203\,
            I => \N__8187\
        );

    \I__1518\ : Span4Mux_v
    port map (
            O => \N__8200\,
            I => \N__8184\
        );

    \I__1517\ : Span4Mux_v
    port map (
            O => \N__8197\,
            I => \N__8181\
        );

    \I__1516\ : InMux
    port map (
            O => \N__8196\,
            I => \N__8176\
        );

    \I__1515\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8176\
        );

    \I__1514\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8169\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8169\
        );

    \I__1512\ : InMux
    port map (
            O => \N__8190\,
            I => \N__8169\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__8187\,
            I => \inst_midgetv_core.INSTR_12\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__8184\,
            I => \inst_midgetv_core.INSTR_12\
        );

    \I__1509\ : Odrv4
    port map (
            O => \N__8181\,
            I => \inst_midgetv_core.INSTR_12\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__8176\,
            I => \inst_midgetv_core.INSTR_12\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__8169\,
            I => \inst_midgetv_core.INSTR_12\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__8158\,
            I => \N__8155\
        );

    \I__1505\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8152\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__8152\,
            I => \inst_midgetv_core.inst_condcode.n5618\
        );

    \I__1503\ : InMux
    port map (
            O => \N__8149\,
            I => \N__8146\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__8146\,
            I => \inst_midgetv_core.inst_ucodepc.n5603\
        );

    \I__1501\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8140\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__8140\,
            I => \inst_midgetv_core.inst_ucodepc.n17\
        );

    \I__1499\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8134\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__8134\,
            I => \inst_midgetv_core.inst_ucodepc.dinx_1_N_145_0\
        );

    \I__1497\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8128\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__8128\,
            I => \N__8125\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__8125\,
            I => \inst_midgetv_core.inst_ucodepc.n5613\
        );

    \I__1494\ : InMux
    port map (
            O => \N__8122\,
            I => \N__8119\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__8119\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk2_illegal_a\
        );

    \I__1492\ : InMux
    port map (
            O => \N__8116\,
            I => \N__8113\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__8113\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n6\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__8110\,
            I => \N__8107\
        );

    \I__1489\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8104\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__8104\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n2\
        );

    \I__1487\ : InMux
    port map (
            O => \N__8101\,
            I => \N__8098\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__8098\,
            I => \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk1_checkfunct7_N_286\
        );

    \I__1485\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8092\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__8092\,
            I => \N__8087\
        );

    \I__1483\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8082\
        );

    \I__1482\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8082\
        );

    \I__1481\ : Sp12to4
    port map (
            O => \N__8087\,
            I => \N__8079\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__8082\,
            I => \N__8076\
        );

    \I__1479\ : Odrv12
    port map (
            O => \N__8079\,
            I => \inst_midgetv_core.ADR_O_28\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__8076\,
            I => \inst_midgetv_core.ADR_O_28\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__8071\,
            I => \inst_midgetv_core.Di_28_cascade_\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__8068\,
            I => \N__8065\
        );

    \I__1475\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8062\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__8062\,
            I => \N__8059\
        );

    \I__1473\ : Sp12to4
    port map (
            O => \N__8059\,
            I => \N__8056\
        );

    \I__1472\ : Odrv12
    port map (
            O => \N__8056\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_28\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__8053\,
            I => \N__8050\
        );

    \I__1470\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8047\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__8047\,
            I => \N__8044\
        );

    \I__1468\ : Span4Mux_h
    port map (
            O => \N__8044\,
            I => \N__8041\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__8041\,
            I => \inst_midgetv_core.rinx_1\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__8038\,
            I => \N__8035\
        );

    \I__1465\ : CascadeBuf
    port map (
            O => \N__8035\,
            I => \N__8032\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__8032\,
            I => \N__8028\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__8031\,
            I => \N__8025\
        );

    \I__1462\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8022\
        );

    \I__1461\ : InMux
    port map (
            O => \N__8025\,
            I => \N__8019\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__8022\,
            I => \N__8016\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__8019\,
            I => \inst_midgetv_core.minx_1\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__8016\,
            I => \inst_midgetv_core.minx_1\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__8011\,
            I => \N__8008\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8008\,
            I => \N__8005\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__8005\,
            I => \N__8002\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__8002\,
            I => \N__7999\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__7999\,
            I => \inst_midgetv_core.rinx_5\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__7996\,
            I => \N__7993\
        );

    \I__1451\ : CascadeBuf
    port map (
            O => \N__7993\,
            I => \N__7990\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__7990\,
            I => \N__7986\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7983\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7980\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7983\,
            I => \N__7977\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7980\,
            I => \N__7974\
        );

    \I__1445\ : Span4Mux_v
    port map (
            O => \N__7977\,
            I => \N__7969\
        );

    \I__1444\ : Span4Mux_h
    port map (
            O => \N__7974\,
            I => \N__7969\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__7969\,
            I => \inst_midgetv_core.minx_5\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__7966\,
            I => \N__7963\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7963\,
            I => \N__7960\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__7960\,
            I => \N__7957\
        );

    \I__1439\ : Span4Mux_h
    port map (
            O => \N__7957\,
            I => \N__7954\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__7954\,
            I => \inst_midgetv_core.rinx_7\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__7951\,
            I => \N__7948\
        );

    \I__1436\ : CascadeBuf
    port map (
            O => \N__7948\,
            I => \N__7944\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7941\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__7944\,
            I => \N__7938\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7941\,
            I => \N__7935\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7932\
        );

    \I__1431\ : Span4Mux_h
    port map (
            O => \N__7935\,
            I => \N__7929\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7932\,
            I => \N__7926\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__7929\,
            I => \inst_midgetv_core.minx_7\
        );

    \I__1428\ : Odrv4
    port map (
            O => \N__7926\,
            I => \inst_midgetv_core.minx_7\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7921\,
            I => \N__7918\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7918\,
            I => \N__7915\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__7915\,
            I => \N__7912\
        );

    \I__1424\ : Odrv4
    port map (
            O => \N__7912\,
            I => \inst_midgetv_core.rinx_3\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__1422\ : CascadeBuf
    port map (
            O => \N__7906\,
            I => \N__7903\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__7903\,
            I => \N__7899\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7896\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7893\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7896\,
            I => \N__7890\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__7893\,
            I => \N__7887\
        );

    \I__1416\ : Odrv4
    port map (
            O => \N__7890\,
            I => \inst_midgetv_core.minx_3\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__7887\,
            I => \inst_midgetv_core.minx_3\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7878\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__7881\,
            I => \N__7870\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7878\,
            I => \N__7866\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7861\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7861\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7850\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7850\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7850\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7870\,
            I => \N__7850\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7850\
        );

    \I__1404\ : Odrv4
    port map (
            O => \N__7866\,
            I => \inst_midgetv_core.inst_ucodepc.usedinx_or_RST_I_notcorerunning\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7861\,
            I => \inst_midgetv_core.inst_ucodepc.usedinx_or_RST_I_notcorerunning\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__7850\,
            I => \inst_midgetv_core.inst_ucodepc.usedinx_or_RST_I_notcorerunning\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__7843\,
            I => \N__7840\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7840\,
            I => \N__7837\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7837\,
            I => \N__7834\
        );

    \I__1398\ : Span4Mux_h
    port map (
            O => \N__7834\,
            I => \N__7831\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__7831\,
            I => \inst_midgetv_core.rinx_6\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7828\,
            I => \N__7810\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7827\,
            I => \N__7810\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7826\,
            I => \N__7810\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7825\,
            I => \N__7810\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7810\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7805\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7805\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7821\,
            I => \N__7802\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__7810\,
            I => \inst_midgetv_core.inst_ucodepc.illegal\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7805\,
            I => \inst_midgetv_core.inst_ucodepc.illegal\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7802\,
            I => \inst_midgetv_core.inst_ucodepc.illegal\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__7795\,
            I => \N__7792\
        );

    \I__1384\ : CascadeBuf
    port map (
            O => \N__7792\,
            I => \N__7789\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__7789\,
            I => \N__7786\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7783\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__7783\,
            I => \N__7780\
        );

    \I__1380\ : Span4Mux_h
    port map (
            O => \N__7780\,
            I => \N__7777\
        );

    \I__1379\ : Odrv4
    port map (
            O => \N__7777\,
            I => \inst_midgetv_core.minx_6\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7774\,
            I => \N__7771\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7771\,
            I => \inst_midgetv_core.inst_ucodepc.n15\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7768\,
            I => \N__7765\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7765\,
            I => \N__7762\
        );

    \I__1374\ : Span4Mux_v
    port map (
            O => \N__7762\,
            I => \N__7759\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__7759\,
            I => \N__7756\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__7756\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09h\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__7753\,
            I => \N__7750\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7745\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7749\,
            I => \N__7740\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7740\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7745\,
            I => \N__7737\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7740\,
            I => \N__7734\
        );

    \I__1365\ : Odrv4
    port map (
            O => \N__7737\,
            I => \inst_midgetv_core.ADR_O_20\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__7734\,
            I => \inst_midgetv_core.ADR_O_20\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__7729\,
            I => \inst_midgetv_core.Di_20_cascade_\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7723\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7723\,
            I => \N__7720\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__7720\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_20\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__7717\,
            I => \N__7714\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7714\,
            I => \N__7711\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7711\,
            I => \N__7708\
        );

    \I__1356\ : Span4Mux_h
    port map (
            O => \N__7708\,
            I => \N__7705\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__7705\,
            I => \N__7702\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__7702\,
            I => \inst_midgetv_core.DAT_O_25\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__7699\,
            I => \inst_midgetv_core.Di_25_cascade_\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__7696\,
            I => \N__7692\
        );

    \I__1351\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7688\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7692\,
            I => \N__7685\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7691\,
            I => \N__7682\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7688\,
            I => \N__7679\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7685\,
            I => \N__7674\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7682\,
            I => \N__7674\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__7679\,
            I => \inst_midgetv_core.ADR_O_25\
        );

    \I__1344\ : Odrv4
    port map (
            O => \N__7674\,
            I => \inst_midgetv_core.ADR_O_25\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7669\,
            I => \N__7666\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7666\,
            I => \N__7663\
        );

    \I__1341\ : Span4Mux_h
    port map (
            O => \N__7663\,
            I => \N__7660\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__7660\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_25\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__7657\,
            I => \N__7654\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7651\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7651\,
            I => \N__7648\
        );

    \I__1336\ : Span4Mux_h
    port map (
            O => \N__7648\,
            I => \N__7645\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__7645\,
            I => \N__7642\
        );

    \I__1334\ : Odrv4
    port map (
            O => \N__7642\,
            I => \inst_midgetv_core.DAT_O_26\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7634\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7638\,
            I => \N__7629\
        );

    \I__1331\ : InMux
    port map (
            O => \N__7637\,
            I => \N__7629\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7634\,
            I => \N__7626\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7629\,
            I => \N__7623\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__7626\,
            I => \inst_midgetv_core.ADR_O_26\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__7623\,
            I => \inst_midgetv_core.ADR_O_26\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__7618\,
            I => \inst_midgetv_core.Di_26_cascade_\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__7615\,
            I => \N__7612\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7609\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__7609\,
            I => \N__7606\
        );

    \I__1322\ : Odrv4
    port map (
            O => \N__7606\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_26\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__7603\,
            I => \N__7600\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7597\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7597\,
            I => \N__7594\
        );

    \I__1318\ : Span4Mux_h
    port map (
            O => \N__7594\,
            I => \N__7591\
        );

    \I__1317\ : Span4Mux_v
    port map (
            O => \N__7591\,
            I => \N__7588\
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__7588\,
            I => \inst_midgetv_core.DAT_O_27\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__7585\,
            I => \N__7582\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7582\,
            I => \N__7577\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7581\,
            I => \N__7572\
        );

    \I__1312\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7572\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7577\,
            I => \N__7569\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__7572\,
            I => \N__7566\
        );

    \I__1309\ : Odrv4
    port map (
            O => \N__7569\,
            I => \inst_midgetv_core.ADR_O_27\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__7566\,
            I => \inst_midgetv_core.ADR_O_27\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__7561\,
            I => \inst_midgetv_core.Di_27_cascade_\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7558\,
            I => \N__7555\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__7555\,
            I => \N__7552\
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__7552\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_27\
        );

    \I__1303\ : InMux
    port map (
            O => \N__7549\,
            I => \N__7546\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__7546\,
            I => \N__7541\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7538\
        );

    \I__1300\ : InMux
    port map (
            O => \N__7544\,
            I => \N__7535\
        );

    \I__1299\ : Span4Mux_h
    port map (
            O => \N__7541\,
            I => \N__7530\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7538\,
            I => \N__7530\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__7535\,
            I => \inst_midgetv_core.ADR_O_29\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__7530\,
            I => \inst_midgetv_core.ADR_O_29\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__7525\,
            I => \N__7522\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7519\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7519\,
            I => \N__7516\
        );

    \I__1292\ : Span4Mux_h
    port map (
            O => \N__7516\,
            I => \N__7513\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__7513\,
            I => \N__7510\
        );

    \I__1290\ : Span4Mux_v
    port map (
            O => \N__7510\,
            I => \N__7507\
        );

    \I__1289\ : Odrv4
    port map (
            O => \N__7507\,
            I => \inst_midgetv_core.DAT_O_28\
        );

    \I__1288\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7501\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__7501\,
            I => \N__7498\
        );

    \I__1286\ : Span4Mux_h
    port map (
            O => \N__7498\,
            I => \N__7495\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__7495\,
            I => \N__7492\
        );

    \I__1284\ : Odrv4
    port map (
            O => \N__7492\,
            I => \inst_midgetv_core.DAT_O_7\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__7489\,
            I => \inst_midgetv_core.Di_7_cascade_\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__7486\,
            I => \N__7483\
        );

    \I__1281\ : InMux
    port map (
            O => \N__7483\,
            I => \N__7480\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__7480\,
            I => \N__7477\
        );

    \I__1279\ : Odrv12
    port map (
            O => \N__7477\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_7\
        );

    \I__1278\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7471\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__7471\,
            I => \N__7468\
        );

    \I__1276\ : Span4Mux_v
    port map (
            O => \N__7468\,
            I => \N__7465\
        );

    \I__1275\ : Span4Mux_h
    port map (
            O => \N__7465\,
            I => \N__7462\
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__7462\,
            I => \inst_midgetv_core.DAT_O_17\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__7459\,
            I => \inst_midgetv_core.Di_17_cascade_\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7453\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__7453\,
            I => \N__7450\
        );

    \I__1270\ : Sp12to4
    port map (
            O => \N__7450\,
            I => \N__7447\
        );

    \I__1269\ : Odrv12
    port map (
            O => \N__7447\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_17\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7441\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__7441\,
            I => \N__7438\
        );

    \I__1266\ : Span4Mux_h
    port map (
            O => \N__7438\,
            I => \N__7435\
        );

    \I__1265\ : Span4Mux_v
    port map (
            O => \N__7435\,
            I => \N__7432\
        );

    \I__1264\ : Odrv4
    port map (
            O => \N__7432\,
            I => \inst_midgetv_core.DAT_O_18\
        );

    \I__1263\ : InMux
    port map (
            O => \N__7429\,
            I => \N__7424\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7428\,
            I => \N__7419\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7419\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__7424\,
            I => \N__7416\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__7419\,
            I => \N__7413\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__7416\,
            I => \inst_midgetv_core.ADR_O_18\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__7413\,
            I => \inst_midgetv_core.ADR_O_18\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__7408\,
            I => \inst_midgetv_core.Di_18_cascade_\
        );

    \I__1255\ : CascadeMux
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__1254\ : InMux
    port map (
            O => \N__7402\,
            I => \N__7399\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__7399\,
            I => \N__7396\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__7396\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_18\
        );

    \I__1251\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7390\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__7390\,
            I => \N__7387\
        );

    \I__1249\ : Span4Mux_h
    port map (
            O => \N__7387\,
            I => \N__7384\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__7384\,
            I => \inst_midgetv_core.DAT_O_19\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__7381\,
            I => \N__7378\
        );

    \I__1246\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7373\
        );

    \I__1245\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7368\
        );

    \I__1244\ : InMux
    port map (
            O => \N__7376\,
            I => \N__7368\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__7373\,
            I => \N__7365\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__7368\,
            I => \N__7362\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__7365\,
            I => \inst_midgetv_core.ADR_O_19\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__7362\,
            I => \inst_midgetv_core.ADR_O_19\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__7357\,
            I => \inst_midgetv_core.Di_19_cascade_\
        );

    \I__1238\ : InMux
    port map (
            O => \N__7354\,
            I => \N__7351\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__7351\,
            I => \N__7348\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__7348\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_19\
        );

    \I__1235\ : InMux
    port map (
            O => \N__7345\,
            I => \N__7342\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__7342\,
            I => \N__7339\
        );

    \I__1233\ : Span4Mux_v
    port map (
            O => \N__7339\,
            I => \N__7336\
        );

    \I__1232\ : Span4Mux_v
    port map (
            O => \N__7336\,
            I => \N__7333\
        );

    \I__1231\ : Odrv4
    port map (
            O => \N__7333\,
            I => \inst_midgetv_core.DAT_O_20\
        );

    \I__1230\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7327\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__7327\,
            I => \N__7322\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7326\,
            I => \N__7319\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7316\
        );

    \I__1226\ : Span4Mux_h
    port map (
            O => \N__7322\,
            I => \N__7309\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__7319\,
            I => \N__7309\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__7316\,
            I => \N__7309\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__7309\,
            I => \inst_midgetv_core.ADR_O_21\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__7306\,
            I => \N__7303\
        );

    \I__1221\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7300\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__7300\,
            I => \N__7297\
        );

    \I__1219\ : Span4Mux_h
    port map (
            O => \N__7297\,
            I => \N__7294\
        );

    \I__1218\ : Span4Mux_v
    port map (
            O => \N__7294\,
            I => \N__7291\
        );

    \I__1217\ : Odrv4
    port map (
            O => \N__7291\,
            I => \inst_midgetv_core.DAT_O_12\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__7288\,
            I => \N__7285\
        );

    \I__1215\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7282\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__7282\,
            I => \N__7277\
        );

    \I__1213\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7272\
        );

    \I__1212\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7272\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__7277\,
            I => \inst_midgetv_core.ADR_O_12\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__7272\,
            I => \inst_midgetv_core.ADR_O_12\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__7267\,
            I => \inst_midgetv_core.Di_12_cascade_\
        );

    \I__1208\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7261\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__7261\,
            I => \N__7258\
        );

    \I__1206\ : Span4Mux_h
    port map (
            O => \N__7258\,
            I => \N__7255\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__7255\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_12\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__7252\,
            I => \N__7249\
        );

    \I__1203\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7246\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__7246\,
            I => \N__7243\
        );

    \I__1201\ : Span4Mux_h
    port map (
            O => \N__7243\,
            I => \N__7240\
        );

    \I__1200\ : Sp12to4
    port map (
            O => \N__7240\,
            I => \N__7237\
        );

    \I__1199\ : Odrv12
    port map (
            O => \N__7237\,
            I => \inst_midgetv_core.DAT_O_29\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__7234\,
            I => \inst_midgetv_core.Di_29_cascade_\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__7231\,
            I => \N__7228\
        );

    \I__1196\ : InMux
    port map (
            O => \N__7228\,
            I => \N__7225\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__7225\,
            I => \N__7222\
        );

    \I__1194\ : Span4Mux_v
    port map (
            O => \N__7222\,
            I => \N__7219\
        );

    \I__1193\ : Odrv4
    port map (
            O => \N__7219\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_29\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__7216\,
            I => \N__7213\
        );

    \I__1191\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7210\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__7210\,
            I => \N__7207\
        );

    \I__1189\ : Span4Mux_v
    port map (
            O => \N__7207\,
            I => \N__7204\
        );

    \I__1188\ : Span4Mux_v
    port map (
            O => \N__7204\,
            I => \N__7201\
        );

    \I__1187\ : Span4Mux_v
    port map (
            O => \N__7201\,
            I => \N__7198\
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__7198\,
            I => \inst_midgetv_core.DAT_O_30\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__7195\,
            I => \N__7192\
        );

    \I__1184\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7189\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__7189\,
            I => \N__7184\
        );

    \I__1182\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7179\
        );

    \I__1181\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7179\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__7184\,
            I => \inst_midgetv_core.ADR_O_30\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__7179\,
            I => \inst_midgetv_core.ADR_O_30\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__7174\,
            I => \inst_midgetv_core.Di_30_cascade_\
        );

    \I__1177\ : InMux
    port map (
            O => \N__7171\,
            I => \N__7168\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__7168\,
            I => \N__7165\
        );

    \I__1175\ : Span4Mux_h
    port map (
            O => \N__7165\,
            I => \N__7162\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__7162\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_30\
        );

    \I__1173\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7156\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__7156\,
            I => \N__7153\
        );

    \I__1171\ : Span4Mux_h
    port map (
            O => \N__7153\,
            I => \N__7150\
        );

    \I__1170\ : Span4Mux_h
    port map (
            O => \N__7150\,
            I => \N__7147\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__7147\,
            I => \inst_midgetv_core.sra_msb\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__7144\,
            I => \N__7139\
        );

    \I__1167\ : InMux
    port map (
            O => \N__7143\,
            I => \N__7132\
        );

    \I__1166\ : InMux
    port map (
            O => \N__7142\,
            I => \N__7132\
        );

    \I__1165\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7132\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__7132\,
            I => \N__7128\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__7131\,
            I => \N__7123\
        );

    \I__1162\ : Span4Mux_h
    port map (
            O => \N__7128\,
            I => \N__7120\
        );

    \I__1161\ : InMux
    port map (
            O => \N__7127\,
            I => \N__7115\
        );

    \I__1160\ : InMux
    port map (
            O => \N__7126\,
            I => \N__7115\
        );

    \I__1159\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7112\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__7120\,
            I => \inst_midgetv_core.ADR_O_31\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__7115\,
            I => \inst_midgetv_core.ADR_O_31\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__7112\,
            I => \inst_midgetv_core.ADR_O_31\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__7105\,
            I => \inst_midgetv_core.Di_31_cascade_\
        );

    \I__1154\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7093\
        );

    \I__1153\ : InMux
    port map (
            O => \N__7101\,
            I => \N__7093\
        );

    \I__1152\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7093\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__7093\,
            I => \N__7090\
        );

    \I__1150\ : Span4Mux_h
    port map (
            O => \N__7090\,
            I => \N__7087\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__7087\,
            I => \inst_midgetv_core.A31\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__7084\,
            I => \inst_midgetv_core.Di_6_cascade_\
        );

    \I__1147\ : InMux
    port map (
            O => \N__7081\,
            I => \N__7078\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__7078\,
            I => \N__7075\
        );

    \I__1145\ : Span4Mux_h
    port map (
            O => \N__7075\,
            I => \N__7072\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__7072\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_6\
        );

    \I__1143\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7066\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__7066\,
            I => \N__7063\
        );

    \I__1141\ : Span4Mux_h
    port map (
            O => \N__7063\,
            I => \N__7060\
        );

    \I__1140\ : Span4Mux_v
    port map (
            O => \N__7060\,
            I => \N__7057\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__7057\,
            I => \inst_midgetv_core.DAT_O_8\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__7054\,
            I => \inst_midgetv_core.Di_8_cascade_\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__7051\,
            I => \N__7048\
        );

    \I__1136\ : InMux
    port map (
            O => \N__7048\,
            I => \N__7045\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__7045\,
            I => \N__7042\
        );

    \I__1134\ : Span4Mux_h
    port map (
            O => \N__7042\,
            I => \N__7039\
        );

    \I__1133\ : Odrv4
    port map (
            O => \N__7039\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_8\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__7036\,
            I => \N__7033\
        );

    \I__1131\ : InMux
    port map (
            O => \N__7033\,
            I => \N__7030\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__7030\,
            I => \N__7027\
        );

    \I__1129\ : Span4Mux_h
    port map (
            O => \N__7027\,
            I => \N__7024\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__7024\,
            I => \inst_midgetv_core.DAT_O_10\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__7021\,
            I => \inst_midgetv_core.Di_10_cascade_\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__7018\,
            I => \N__7015\
        );

    \I__1125\ : InMux
    port map (
            O => \N__7015\,
            I => \N__7012\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__7012\,
            I => \N__7009\
        );

    \I__1123\ : Span4Mux_h
    port map (
            O => \N__7009\,
            I => \N__7006\
        );

    \I__1122\ : Odrv4
    port map (
            O => \N__7006\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_10\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__7003\,
            I => \N__7000\
        );

    \I__1120\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6997\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6997\,
            I => \N__6994\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__6994\,
            I => \N__6991\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__6991\,
            I => \inst_midgetv_core.DAT_O_11\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__6988\,
            I => \inst_midgetv_core.Di_11_cascade_\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6985\,
            I => \N__6982\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__1113\ : Span4Mux_h
    port map (
            O => \N__6979\,
            I => \N__6976\
        );

    \I__1112\ : Odrv4
    port map (
            O => \N__6976\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_11\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6973\,
            I => \N__6970\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6970\,
            I => \N__6966\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6969\,
            I => \N__6963\
        );

    \I__1108\ : Span4Mux_h
    port map (
            O => \N__6966\,
            I => \N__6958\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6963\,
            I => \N__6955\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6950\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6950\
        );

    \I__1104\ : Odrv4
    port map (
            O => \N__6958\,
            I => \inst_midgetv_core.ADR_O_10\
        );

    \I__1103\ : Odrv4
    port map (
            O => \N__6955\,
            I => \inst_midgetv_core.ADR_O_10\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6950\,
            I => \inst_midgetv_core.ADR_O_10\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__6943\,
            I => \N__6940\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6937\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6937\,
            I => \N__6934\
        );

    \I__1098\ : Span4Mux_h
    port map (
            O => \N__6934\,
            I => \N__6931\
        );

    \I__1097\ : Odrv4
    port map (
            O => \N__6931\,
            I => \inst_midgetv_core.DAT_O_9\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__6928\,
            I => \inst_midgetv_core.Di_9_cascade_\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6921\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6918\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6921\,
            I => \N__6915\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6918\,
            I => \N__6910\
        );

    \I__1091\ : Span4Mux_h
    port map (
            O => \N__6915\,
            I => \N__6907\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6914\,
            I => \N__6904\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6901\
        );

    \I__1088\ : Odrv12
    port map (
            O => \N__6910\,
            I => \inst_midgetv_core.ADR_O_9\
        );

    \I__1087\ : Odrv4
    port map (
            O => \N__6907\,
            I => \inst_midgetv_core.ADR_O_9\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6904\,
            I => \inst_midgetv_core.ADR_O_9\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6901\,
            I => \inst_midgetv_core.ADR_O_9\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__6892\,
            I => \N__6889\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6889\,
            I => \N__6886\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__6886\,
            I => \N__6883\
        );

    \I__1081\ : Span4Mux_v
    port map (
            O => \N__6883\,
            I => \N__6880\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__6880\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_9\
        );

    \I__1079\ : CascadeMux
    port map (
            O => \N__6877\,
            I => \inst_midgetv_core.Di_2_cascade_\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6874\,
            I => \N__6871\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6871\,
            I => \N__6868\
        );

    \I__1076\ : Span4Mux_h
    port map (
            O => \N__6868\,
            I => \N__6865\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__6865\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_2\
        );

    \I__1074\ : CascadeMux
    port map (
            O => \N__6862\,
            I => \N__6858\
        );

    \I__1073\ : IoInMux
    port map (
            O => \N__6861\,
            I => \N__6855\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6852\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6855\,
            I => \N__6849\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6852\,
            I => \N__6846\
        );

    \I__1069\ : Span12Mux_s5_v
    port map (
            O => \N__6849\,
            I => \N__6843\
        );

    \I__1068\ : Span4Mux_h
    port map (
            O => \N__6846\,
            I => \N__6840\
        );

    \I__1067\ : Odrv12
    port map (
            O => \N__6843\,
            I => \DAT_O_3\
        );

    \I__1066\ : Odrv4
    port map (
            O => \N__6840\,
            I => \DAT_O_3\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__6835\,
            I => \inst_midgetv_core.Di_3_cascade_\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6832\,
            I => \N__6829\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6829\,
            I => \N__6826\
        );

    \I__1062\ : Span4Mux_h
    port map (
            O => \N__6826\,
            I => \N__6823\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__6823\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_3\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__6820\,
            I => \N__6817\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6817\,
            I => \N__6814\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6814\,
            I => \N__6811\
        );

    \I__1057\ : Span4Mux_h
    port map (
            O => \N__6811\,
            I => \N__6808\
        );

    \I__1056\ : Odrv4
    port map (
            O => \N__6808\,
            I => \inst_midgetv_core.DAT_O_4\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__6805\,
            I => \inst_midgetv_core.Di_4_cascade_\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6802\,
            I => \N__6799\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6799\,
            I => \N__6796\
        );

    \I__1052\ : Span4Mux_h
    port map (
            O => \N__6796\,
            I => \N__6793\
        );

    \I__1051\ : Odrv4
    port map (
            O => \N__6793\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_4\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6787\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6787\,
            I => \N__6784\
        );

    \I__1048\ : Span4Mux_v
    port map (
            O => \N__6784\,
            I => \N__6781\
        );

    \I__1047\ : Odrv4
    port map (
            O => \N__6781\,
            I => \inst_midgetv_core.DAT_O_5\
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__6778\,
            I => \inst_midgetv_core.Di_5_cascade_\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6772\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6772\,
            I => \N__6769\
        );

    \I__1043\ : Span4Mux_v
    port map (
            O => \N__6769\,
            I => \N__6766\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__6766\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_5\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__6763\,
            I => \N__6760\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6760\,
            I => \N__6757\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6757\,
            I => \N__6754\
        );

    \I__1038\ : Span4Mux_h
    port map (
            O => \N__6754\,
            I => \N__6751\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__6751\,
            I => \inst_midgetv_core.DAT_O_6\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6745\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6745\,
            I => \N__6742\
        );

    \I__1034\ : Span4Mux_v
    port map (
            O => \N__6742\,
            I => \N__6739\
        );

    \I__1033\ : Odrv4
    port map (
            O => \N__6739\,
            I => \inst_midgetv_core.sa43\
        );

    \I__1032\ : CEMux
    port map (
            O => \N__6736\,
            I => \N__6733\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6733\,
            I => \N__6730\
        );

    \I__1030\ : Span4Mux_v
    port map (
            O => \N__6730\,
            I => \N__6727\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__6727\,
            I => \N__6724\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__6724\,
            I => \inst_midgetv_core.inst_progressctrl.n2764\
        );

    \I__1027\ : SRMux
    port map (
            O => \N__6721\,
            I => \N__6718\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6718\,
            I => \N__6715\
        );

    \I__1025\ : Span4Mux_h
    port map (
            O => \N__6715\,
            I => \N__6712\
        );

    \I__1024\ : Span4Mux_v
    port map (
            O => \N__6712\,
            I => \N__6709\
        );

    \I__1023\ : Span4Mux_h
    port map (
            O => \N__6709\,
            I => \N__6705\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6708\,
            I => \N__6702\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__6705\,
            I => \inst_midgetv_core.inst_progressctrl.ctrlreg_we_N_84\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6702\,
            I => \inst_midgetv_core.inst_progressctrl.ctrlreg_we_N_84\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6691\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6691\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6691\,
            I => \N__6688\
        );

    \I__1016\ : Span4Mux_h
    port map (
            O => \N__6688\,
            I => \N__6685\
        );

    \I__1015\ : Odrv4
    port map (
            O => \N__6685\,
            I => \inst_midgetv_core.sa14\
        );

    \I__1014\ : SRMux
    port map (
            O => \N__6682\,
            I => \N__6675\
        );

    \I__1013\ : SRMux
    port map (
            O => \N__6681\,
            I => \N__6672\
        );

    \I__1012\ : SRMux
    port map (
            O => \N__6680\,
            I => \N__6669\
        );

    \I__1011\ : SRMux
    port map (
            O => \N__6679\,
            I => \N__6666\
        );

    \I__1010\ : SRMux
    port map (
            O => \N__6678\,
            I => \N__6663\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6675\,
            I => \N__6660\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6672\,
            I => \N__6655\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6669\,
            I => \N__6655\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6666\,
            I => \N__6652\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__6663\,
            I => \N__6649\
        );

    \I__1004\ : Span4Mux_v
    port map (
            O => \N__6660\,
            I => \N__6646\
        );

    \I__1003\ : Span4Mux_v
    port map (
            O => \N__6655\,
            I => \N__6639\
        );

    \I__1002\ : Span4Mux_v
    port map (
            O => \N__6652\,
            I => \N__6639\
        );

    \I__1001\ : Span4Mux_h
    port map (
            O => \N__6649\,
            I => \N__6639\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__6646\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_nsa14_or_nCORERUNNING\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__6639\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_nsa14_or_nCORERUNNING\
        );

    \I__998\ : IoInMux
    port map (
            O => \N__6634\,
            I => \N__6630\
        );

    \I__997\ : IoInMux
    port map (
            O => \N__6633\,
            I => \N__6627\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__6630\,
            I => \N__6624\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6627\,
            I => \N__6621\
        );

    \I__994\ : IoSpan4Mux
    port map (
            O => \N__6624\,
            I => \N__6618\
        );

    \I__993\ : IoSpan4Mux
    port map (
            O => \N__6621\,
            I => \N__6614\
        );

    \I__992\ : Span4Mux_s3_v
    port map (
            O => \N__6618\,
            I => \N__6611\
        );

    \I__991\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6608\
        );

    \I__990\ : Sp12to4
    port map (
            O => \N__6614\,
            I => \N__6605\
        );

    \I__989\ : Span4Mux_v
    port map (
            O => \N__6611\,
            I => \N__6602\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6608\,
            I => \N__6599\
        );

    \I__987\ : Span12Mux_s9_v
    port map (
            O => \N__6605\,
            I => \N__6596\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__6602\,
            I => \N__6591\
        );

    \I__985\ : Span4Mux_h
    port map (
            O => \N__6599\,
            I => \N__6591\
        );

    \I__984\ : Odrv12
    port map (
            O => \N__6596\,
            I => \DAT_O_0\
        );

    \I__983\ : Odrv4
    port map (
            O => \N__6591\,
            I => \DAT_O_0\
        );

    \I__982\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6583\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__6583\,
            I => \inst_midgetv_core.INSTR_0\
        );

    \I__980\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6576\
        );

    \I__979\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6573\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6576\,
            I => \inst_midgetv_core.ADR_O_0\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__6573\,
            I => \inst_midgetv_core.ADR_O_0\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__6568\,
            I => \inst_midgetv_core.Di_0_cascade_\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__6565\,
            I => \N__6562\
        );

    \I__974\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6559\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__972\ : Span4Mux_h
    port map (
            O => \N__6556\,
            I => \N__6553\
        );

    \I__971\ : Odrv4
    port map (
            O => \N__6553\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_0\
        );

    \I__970\ : IoInMux
    port map (
            O => \N__6550\,
            I => \N__6547\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6547\,
            I => \N__6544\
        );

    \I__968\ : Span4Mux_s2_v
    port map (
            O => \N__6544\,
            I => \N__6541\
        );

    \I__967\ : Span4Mux_v
    port map (
            O => \N__6541\,
            I => \N__6537\
        );

    \I__966\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6534\
        );

    \I__965\ : Span4Mux_v
    port map (
            O => \N__6537\,
            I => \N__6531\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__6534\,
            I => \N__6528\
        );

    \I__963\ : Span4Mux_v
    port map (
            O => \N__6531\,
            I => \N__6525\
        );

    \I__962\ : Span4Mux_h
    port map (
            O => \N__6528\,
            I => \N__6522\
        );

    \I__961\ : Odrv4
    port map (
            O => \N__6525\,
            I => \DAT_O_1\
        );

    \I__960\ : Odrv4
    port map (
            O => \N__6522\,
            I => \DAT_O_1\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__6517\,
            I => \N__6514\
        );

    \I__958\ : InMux
    port map (
            O => \N__6514\,
            I => \N__6511\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__6511\,
            I => \inst_midgetv_core.INSTR_1\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__6508\,
            I => \inst_midgetv_core.Di_1_cascade_\
        );

    \I__955\ : CascadeMux
    port map (
            O => \N__6505\,
            I => \N__6500\
        );

    \I__954\ : InMux
    port map (
            O => \N__6504\,
            I => \N__6497\
        );

    \I__953\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6492\
        );

    \I__952\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6492\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__6497\,
            I => \inst_midgetv_core.ADR_O_1\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__6492\,
            I => \inst_midgetv_core.ADR_O_1\
        );

    \I__949\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6484\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__6484\,
            I => \N__6481\
        );

    \I__947\ : Span4Mux_v
    port map (
            O => \N__6481\,
            I => \N__6478\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__6478\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_1\
        );

    \I__945\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6472\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__6472\,
            I => \N__6467\
        );

    \I__943\ : InMux
    port map (
            O => \N__6471\,
            I => \N__6462\
        );

    \I__942\ : InMux
    port map (
            O => \N__6470\,
            I => \N__6462\
        );

    \I__941\ : Span4Mux_h
    port map (
            O => \N__6467\,
            I => \N__6457\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__6462\,
            I => \N__6457\
        );

    \I__939\ : Odrv4
    port map (
            O => \N__6457\,
            I => \inst_midgetv_core.ADR_O_23\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__6454\,
            I => \inst_midgetv_core.Di_23_cascade_\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__6451\,
            I => \N__6448\
        );

    \I__936\ : InMux
    port map (
            O => \N__6448\,
            I => \N__6445\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__6445\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_23\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__6442\,
            I => \N__6439\
        );

    \I__933\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6436\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__6436\,
            I => \N__6433\
        );

    \I__931\ : Span4Mux_h
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__930\ : Span4Mux_v
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__6427\,
            I => \N__6424\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__6424\,
            I => \inst_midgetv_core.DAT_O_24\
        );

    \I__927\ : InMux
    port map (
            O => \N__6421\,
            I => \N__6416\
        );

    \I__926\ : InMux
    port map (
            O => \N__6420\,
            I => \N__6411\
        );

    \I__925\ : InMux
    port map (
            O => \N__6419\,
            I => \N__6411\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__6416\,
            I => \N__6406\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__6411\,
            I => \N__6406\
        );

    \I__922\ : Span4Mux_v
    port map (
            O => \N__6406\,
            I => \N__6403\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__6403\,
            I => \inst_midgetv_core.ADR_O_24\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__6400\,
            I => \inst_midgetv_core.Di_24_cascade_\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__6397\,
            I => \N__6394\
        );

    \I__918\ : InMux
    port map (
            O => \N__6394\,
            I => \N__6391\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6391\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_24\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__6388\,
            I => \N__6385\
        );

    \I__915\ : CascadeBuf
    port map (
            O => \N__6385\,
            I => \N__6382\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__6382\,
            I => \N__6379\
        );

    \I__913\ : CascadeBuf
    port map (
            O => \N__6379\,
            I => \N__6376\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__6376\,
            I => \N__6373\
        );

    \I__911\ : CascadeBuf
    port map (
            O => \N__6373\,
            I => \N__6370\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__6370\,
            I => \N__6367\
        );

    \I__909\ : CascadeBuf
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__6364\,
            I => \N__6361\
        );

    \I__907\ : CascadeBuf
    port map (
            O => \N__6361\,
            I => \N__6358\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__6358\,
            I => \N__6355\
        );

    \I__905\ : CascadeBuf
    port map (
            O => \N__6355\,
            I => \N__6352\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__6352\,
            I => \N__6349\
        );

    \I__903\ : CascadeBuf
    port map (
            O => \N__6349\,
            I => \N__6346\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__6346\,
            I => \N__6343\
        );

    \I__901\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6340\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__6340\,
            I => \N__6337\
        );

    \I__899\ : Span4Mux_s2_v
    port map (
            O => \N__6337\,
            I => \N__6334\
        );

    \I__898\ : Span4Mux_h
    port map (
            O => \N__6334\,
            I => \N__6331\
        );

    \I__897\ : Span4Mux_v
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__6328\,
            I => \inst_midgetv_core.Wai_7\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__6325\,
            I => \N__6322\
        );

    \I__894\ : CascadeBuf
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__892\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__6313\,
            I => \N__6309\
        );

    \I__890\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6306\
        );

    \I__889\ : Span4Mux_h
    port map (
            O => \N__6309\,
            I => \N__6303\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__6306\,
            I => \inst_midgetv_core.mostofminx0\
        );

    \I__887\ : Odrv4
    port map (
            O => \N__6303\,
            I => \inst_midgetv_core.mostofminx0\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__6298\,
            I => \N__6295\
        );

    \I__885\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6292\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__883\ : Span4Mux_h
    port map (
            O => \N__6289\,
            I => \N__6286\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__6286\,
            I => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.instr0100\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__6283\,
            I => \N__6280\
        );

    \I__880\ : InMux
    port map (
            O => \N__6280\,
            I => \N__6277\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__6277\,
            I => \N__6274\
        );

    \I__878\ : Span4Mux_h
    port map (
            O => \N__6274\,
            I => \N__6271\
        );

    \I__877\ : Odrv4
    port map (
            O => \N__6271\,
            I => \inst_midgetv_core.rinx_4\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__6268\,
            I => \N__6265\
        );

    \I__875\ : CascadeBuf
    port map (
            O => \N__6265\,
            I => \N__6262\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__6262\,
            I => \N__6258\
        );

    \I__873\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6255\
        );

    \I__872\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6252\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__6255\,
            I => \N__6249\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__6252\,
            I => \N__6246\
        );

    \I__869\ : Odrv4
    port map (
            O => \N__6249\,
            I => \inst_midgetv_core.minx_4\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__6246\,
            I => \inst_midgetv_core.minx_4\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__6241\,
            I => \N__6238\
        );

    \I__866\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6235\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__6235\,
            I => \N__6232\
        );

    \I__864\ : Span4Mux_v
    port map (
            O => \N__6232\,
            I => \N__6229\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__6229\,
            I => \inst_midgetv_core.rinx_2\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__6226\,
            I => \N__6223\
        );

    \I__861\ : CascadeBuf
    port map (
            O => \N__6223\,
            I => \N__6220\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__6220\,
            I => \N__6217\
        );

    \I__859\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6213\
        );

    \I__858\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6210\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__6213\,
            I => \N__6207\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__6210\,
            I => \inst_midgetv_core.minx_2\
        );

    \I__855\ : Odrv12
    port map (
            O => \N__6207\,
            I => \inst_midgetv_core.minx_2\
        );

    \I__854\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6199\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__6199\,
            I => \N__6196\
        );

    \I__852\ : Span4Mux_h
    port map (
            O => \N__6196\,
            I => \N__6193\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__6193\,
            I => \N__6189\
        );

    \I__850\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6186\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__6189\,
            I => \N__6183\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__6186\,
            I => \N__6180\
        );

    \I__847\ : Span4Mux_v
    port map (
            O => \N__6183\,
            I => \N__6175\
        );

    \I__846\ : Span4Mux_h
    port map (
            O => \N__6180\,
            I => \N__6175\
        );

    \I__845\ : Odrv4
    port map (
            O => \N__6175\,
            I => \inst_midgetv_core.B_29\
        );

    \I__844\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6162\
        );

    \I__843\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6147\
        );

    \I__842\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6147\
        );

    \I__841\ : InMux
    port map (
            O => \N__6169\,
            I => \N__6147\
        );

    \I__840\ : InMux
    port map (
            O => \N__6168\,
            I => \N__6147\
        );

    \I__839\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6147\
        );

    \I__838\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6147\
        );

    \I__837\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6147\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__6162\,
            I => \N__6138\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__6147\,
            I => \N__6138\
        );

    \I__834\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6129\
        );

    \I__833\ : InMux
    port map (
            O => \N__6145\,
            I => \N__6129\
        );

    \I__832\ : InMux
    port map (
            O => \N__6144\,
            I => \N__6129\
        );

    \I__831\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6129\
        );

    \I__830\ : Span4Mux_h
    port map (
            O => \N__6138\,
            I => \N__6126\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__6129\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa13\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__6126\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa13\
        );

    \I__827\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6112\
        );

    \I__826\ : InMux
    port map (
            O => \N__6120\,
            I => \N__6112\
        );

    \I__825\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6112\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__6112\,
            I => \N__6109\
        );

    \I__823\ : Span4Mux_v
    port map (
            O => \N__6109\,
            I => \N__6106\
        );

    \I__822\ : Span4Mux_v
    port map (
            O => \N__6106\,
            I => \N__6103\
        );

    \I__821\ : Span4Mux_v
    port map (
            O => \N__6103\,
            I => \N__6100\
        );

    \I__820\ : Span4Mux_v
    port map (
            O => \N__6100\,
            I => \N__6097\
        );

    \I__819\ : IoSpan4Mux
    port map (
            O => \N__6097\,
            I => \N__6094\
        );

    \I__818\ : Span4Mux_s3_v
    port map (
            O => \N__6094\,
            I => \N__6085\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__6093\,
            I => \N__6082\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__6092\,
            I => \N__6079\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__6091\,
            I => \N__6075\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__6090\,
            I => \N__6072\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__6089\,
            I => \N__6069\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__6088\,
            I => \N__6066\
        );

    \I__811\ : Span4Mux_v
    port map (
            O => \N__6085\,
            I => \N__6058\
        );

    \I__810\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6046\
        );

    \I__809\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6046\
        );

    \I__808\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6046\
        );

    \I__807\ : InMux
    port map (
            O => \N__6075\,
            I => \N__6046\
        );

    \I__806\ : InMux
    port map (
            O => \N__6072\,
            I => \N__6037\
        );

    \I__805\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6037\
        );

    \I__804\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6037\
        );

    \I__803\ : InMux
    port map (
            O => \N__6065\,
            I => \N__6037\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__6064\,
            I => \N__6034\
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__6063\,
            I => \N__6031\
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__6062\,
            I => \N__6028\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__6061\,
            I => \N__6025\
        );

    \I__798\ : Span4Mux_v
    port map (
            O => \N__6058\,
            I => \N__6022\
        );

    \I__797\ : InMux
    port map (
            O => \N__6057\,
            I => \N__6015\
        );

    \I__796\ : InMux
    port map (
            O => \N__6056\,
            I => \N__6015\
        );

    \I__795\ : InMux
    port map (
            O => \N__6055\,
            I => \N__6015\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__6046\,
            I => \N__6010\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__6037\,
            I => \N__6010\
        );

    \I__792\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6005\
        );

    \I__791\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6005\
        );

    \I__790\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6000\
        );

    \I__789\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6000\
        );

    \I__788\ : Span4Mux_v
    port map (
            O => \N__6022\,
            I => \N__5997\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__6015\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa10\
        );

    \I__786\ : Odrv4
    port map (
            O => \N__6010\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa10\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__6005\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa10\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__6000\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa10\
        );

    \I__783\ : Odrv4
    port map (
            O => \N__5997\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa10\
        );

    \I__782\ : InMux
    port map (
            O => \N__5986\,
            I => \bfn_14_19_0_\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__5983\,
            I => \N__5980\
        );

    \I__780\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5977\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5977\,
            I => \N__5974\
        );

    \I__778\ : Span4Mux_v
    port map (
            O => \N__5974\,
            I => \N__5971\
        );

    \I__777\ : Span4Mux_h
    port map (
            O => \N__5971\,
            I => \N__5968\
        );

    \I__776\ : Odrv4
    port map (
            O => \N__5968\,
            I => \inst_midgetv_core.DAT_O_21\
        );

    \I__775\ : CascadeMux
    port map (
            O => \N__5965\,
            I => \inst_midgetv_core.Di_21_cascade_\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__5962\,
            I => \N__5959\
        );

    \I__773\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5956\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5956\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_21\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__5953\,
            I => \N__5950\
        );

    \I__770\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5947\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5947\,
            I => \N__5944\
        );

    \I__768\ : Span4Mux_v
    port map (
            O => \N__5944\,
            I => \N__5941\
        );

    \I__767\ : Span4Mux_h
    port map (
            O => \N__5941\,
            I => \N__5938\
        );

    \I__766\ : Odrv4
    port map (
            O => \N__5938\,
            I => \inst_midgetv_core.DAT_O_22\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__5935\,
            I => \N__5932\
        );

    \I__764\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5927\
        );

    \I__763\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5922\
        );

    \I__762\ : InMux
    port map (
            O => \N__5930\,
            I => \N__5922\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5927\,
            I => \N__5917\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5922\,
            I => \N__5917\
        );

    \I__759\ : Odrv4
    port map (
            O => \N__5917\,
            I => \inst_midgetv_core.ADR_O_22\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__5914\,
            I => \inst_midgetv_core.Di_22_cascade_\
        );

    \I__757\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5908\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5908\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.A_22\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__5905\,
            I => \N__5902\
        );

    \I__754\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5899\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5899\,
            I => \N__5896\
        );

    \I__752\ : Span4Mux_v
    port map (
            O => \N__5896\,
            I => \N__5893\
        );

    \I__751\ : Span4Mux_h
    port map (
            O => \N__5893\,
            I => \N__5890\
        );

    \I__750\ : Odrv4
    port map (
            O => \N__5890\,
            I => \inst_midgetv_core.DAT_O_23\
        );

    \I__749\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5884\,
            I => \N__5880\
        );

    \I__747\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5877\
        );

    \I__746\ : Span4Mux_h
    port map (
            O => \N__5880\,
            I => \N__5874\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5877\,
            I => \N__5871\
        );

    \I__744\ : Span4Mux_h
    port map (
            O => \N__5874\,
            I => \N__5868\
        );

    \I__743\ : Span4Mux_h
    port map (
            O => \N__5871\,
            I => \N__5865\
        );

    \I__742\ : Span4Mux_v
    port map (
            O => \N__5868\,
            I => \N__5862\
        );

    \I__741\ : Span4Mux_h
    port map (
            O => \N__5865\,
            I => \N__5859\
        );

    \I__740\ : Odrv4
    port map (
            O => \N__5862\,
            I => \inst_midgetv_core.B_21\
        );

    \I__739\ : Odrv4
    port map (
            O => \N__5859\,
            I => \inst_midgetv_core.B_21\
        );

    \I__738\ : InMux
    port map (
            O => \N__5854\,
            I => \N__5851\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__5851\,
            I => \N__5848\
        );

    \I__736\ : Span4Mux_h
    port map (
            O => \N__5848\,
            I => \N__5844\
        );

    \I__735\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5841\
        );

    \I__734\ : Span4Mux_h
    port map (
            O => \N__5844\,
            I => \N__5838\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5841\,
            I => \N__5835\
        );

    \I__732\ : Span4Mux_v
    port map (
            O => \N__5838\,
            I => \N__5830\
        );

    \I__731\ : Span4Mux_h
    port map (
            O => \N__5835\,
            I => \N__5830\
        );

    \I__730\ : Odrv4
    port map (
            O => \N__5830\,
            I => \inst_midgetv_core.B_22\
        );

    \I__729\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5824\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__5824\,
            I => \N__5821\
        );

    \I__727\ : Span4Mux_h
    port map (
            O => \N__5821\,
            I => \N__5817\
        );

    \I__726\ : InMux
    port map (
            O => \N__5820\,
            I => \N__5814\
        );

    \I__725\ : Span4Mux_h
    port map (
            O => \N__5817\,
            I => \N__5811\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5814\,
            I => \N__5808\
        );

    \I__723\ : Span4Mux_v
    port map (
            O => \N__5811\,
            I => \N__5805\
        );

    \I__722\ : Span4Mux_v
    port map (
            O => \N__5808\,
            I => \N__5802\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__5805\,
            I => \inst_midgetv_core.B_23\
        );

    \I__720\ : Odrv4
    port map (
            O => \N__5802\,
            I => \inst_midgetv_core.B_23\
        );

    \I__719\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5793\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__5796\,
            I => \N__5790\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5793\,
            I => \N__5787\
        );

    \I__716\ : InMux
    port map (
            O => \N__5790\,
            I => \N__5784\
        );

    \I__715\ : Span4Mux_h
    port map (
            O => \N__5787\,
            I => \N__5781\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5784\,
            I => \N__5778\
        );

    \I__713\ : Span4Mux_v
    port map (
            O => \N__5781\,
            I => \N__5775\
        );

    \I__712\ : Span4Mux_h
    port map (
            O => \N__5778\,
            I => \N__5772\
        );

    \I__711\ : Span4Mux_v
    port map (
            O => \N__5775\,
            I => \N__5769\
        );

    \I__710\ : Sp12to4
    port map (
            O => \N__5772\,
            I => \N__5766\
        );

    \I__709\ : Odrv4
    port map (
            O => \N__5769\,
            I => \inst_midgetv_core.B_24\
        );

    \I__708\ : Odrv12
    port map (
            O => \N__5766\,
            I => \inst_midgetv_core.B_24\
        );

    \I__707\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5758\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5758\,
            I => \N__5755\
        );

    \I__705\ : Span4Mux_v
    port map (
            O => \N__5755\,
            I => \N__5751\
        );

    \I__704\ : InMux
    port map (
            O => \N__5754\,
            I => \N__5748\
        );

    \I__703\ : Span4Mux_h
    port map (
            O => \N__5751\,
            I => \N__5745\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5748\,
            I => \N__5742\
        );

    \I__701\ : Span4Mux_v
    port map (
            O => \N__5745\,
            I => \N__5739\
        );

    \I__700\ : Span4Mux_h
    port map (
            O => \N__5742\,
            I => \N__5736\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__5739\,
            I => \inst_midgetv_core.B_25\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__5736\,
            I => \inst_midgetv_core.B_25\
        );

    \I__697\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5728\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__695\ : Span4Mux_h
    port map (
            O => \N__5725\,
            I => \N__5721\
        );

    \I__694\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5718\
        );

    \I__693\ : Span4Mux_h
    port map (
            O => \N__5721\,
            I => \N__5715\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5718\,
            I => \N__5712\
        );

    \I__691\ : Span4Mux_v
    port map (
            O => \N__5715\,
            I => \N__5709\
        );

    \I__690\ : Span4Mux_h
    port map (
            O => \N__5712\,
            I => \N__5706\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__5709\,
            I => \inst_midgetv_core.B_26\
        );

    \I__688\ : Odrv4
    port map (
            O => \N__5706\,
            I => \inst_midgetv_core.B_26\
        );

    \I__687\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5698\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5698\,
            I => \N__5695\
        );

    \I__685\ : Span4Mux_h
    port map (
            O => \N__5695\,
            I => \N__5691\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__5694\,
            I => \N__5688\
        );

    \I__683\ : Span4Mux_h
    port map (
            O => \N__5691\,
            I => \N__5685\
        );

    \I__682\ : InMux
    port map (
            O => \N__5688\,
            I => \N__5682\
        );

    \I__681\ : Span4Mux_v
    port map (
            O => \N__5685\,
            I => \N__5679\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5682\,
            I => \N__5676\
        );

    \I__679\ : Odrv4
    port map (
            O => \N__5679\,
            I => \inst_midgetv_core.B_27\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__5676\,
            I => \inst_midgetv_core.B_27\
        );

    \I__677\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5668\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5668\,
            I => \N__5665\
        );

    \I__675\ : Span4Mux_h
    port map (
            O => \N__5665\,
            I => \N__5662\
        );

    \I__674\ : Span4Mux_h
    port map (
            O => \N__5662\,
            I => \N__5658\
        );

    \I__673\ : InMux
    port map (
            O => \N__5661\,
            I => \N__5655\
        );

    \I__672\ : Span4Mux_v
    port map (
            O => \N__5658\,
            I => \N__5652\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__5655\,
            I => \N__5649\
        );

    \I__670\ : Span4Mux_v
    port map (
            O => \N__5652\,
            I => \N__5644\
        );

    \I__669\ : Span4Mux_h
    port map (
            O => \N__5649\,
            I => \N__5644\
        );

    \I__668\ : Odrv4
    port map (
            O => \N__5644\,
            I => \inst_midgetv_core.B_28\
        );

    \I__667\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5638\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5638\,
            I => \N__5634\
        );

    \I__665\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5631\
        );

    \I__664\ : Span4Mux_v
    port map (
            O => \N__5634\,
            I => \N__5628\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__5631\,
            I => \N__5625\
        );

    \I__662\ : Span4Mux_h
    port map (
            O => \N__5628\,
            I => \N__5622\
        );

    \I__661\ : Span4Mux_h
    port map (
            O => \N__5625\,
            I => \N__5619\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__5622\,
            I => \inst_midgetv_core.B_13\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__5619\,
            I => \inst_midgetv_core.B_13\
        );

    \I__658\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5611\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5611\,
            I => \N__5607\
        );

    \I__656\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5604\
        );

    \I__655\ : Span4Mux_v
    port map (
            O => \N__5607\,
            I => \N__5601\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__5604\,
            I => \N__5598\
        );

    \I__653\ : Span4Mux_h
    port map (
            O => \N__5601\,
            I => \N__5595\
        );

    \I__652\ : Span4Mux_h
    port map (
            O => \N__5598\,
            I => \N__5592\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__5595\,
            I => \inst_midgetv_core.B_14\
        );

    \I__650\ : Odrv4
    port map (
            O => \N__5592\,
            I => \inst_midgetv_core.B_14\
        );

    \I__649\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5583\
        );

    \I__648\ : InMux
    port map (
            O => \N__5586\,
            I => \N__5580\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__5583\,
            I => \N__5577\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__5580\,
            I => \N__5574\
        );

    \I__645\ : Span12Mux_h
    port map (
            O => \N__5577\,
            I => \N__5571\
        );

    \I__644\ : Span4Mux_h
    port map (
            O => \N__5574\,
            I => \N__5568\
        );

    \I__643\ : Odrv12
    port map (
            O => \N__5571\,
            I => \inst_midgetv_core.B_15\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__5568\,
            I => \inst_midgetv_core.B_15\
        );

    \I__641\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5560\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__5560\,
            I => \N__5557\
        );

    \I__639\ : Span4Mux_h
    port map (
            O => \N__5557\,
            I => \N__5553\
        );

    \I__638\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5550\
        );

    \I__637\ : Span4Mux_h
    port map (
            O => \N__5553\,
            I => \N__5547\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5550\,
            I => \N__5544\
        );

    \I__635\ : Span4Mux_v
    port map (
            O => \N__5547\,
            I => \N__5541\
        );

    \I__634\ : Span4Mux_v
    port map (
            O => \N__5544\,
            I => \N__5538\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__5541\,
            I => \inst_midgetv_core.B_16\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__5538\,
            I => \inst_midgetv_core.B_16\
        );

    \I__631\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5530\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__629\ : Span4Mux_v
    port map (
            O => \N__5527\,
            I => \N__5523\
        );

    \I__628\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5520\
        );

    \I__627\ : Span4Mux_h
    port map (
            O => \N__5523\,
            I => \N__5517\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__5520\,
            I => \N__5514\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__5517\,
            I => \N__5511\
        );

    \I__624\ : Span4Mux_h
    port map (
            O => \N__5514\,
            I => \N__5508\
        );

    \I__623\ : Odrv4
    port map (
            O => \N__5511\,
            I => \inst_midgetv_core.B_17\
        );

    \I__622\ : Odrv4
    port map (
            O => \N__5508\,
            I => \inst_midgetv_core.B_17\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__5503\,
            I => \N__5500\
        );

    \I__620\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5496\
        );

    \I__619\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5493\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__5496\,
            I => \N__5490\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5493\,
            I => \N__5487\
        );

    \I__616\ : Span4Mux_v
    port map (
            O => \N__5490\,
            I => \N__5484\
        );

    \I__615\ : Span4Mux_v
    port map (
            O => \N__5487\,
            I => \N__5479\
        );

    \I__614\ : Span4Mux_h
    port map (
            O => \N__5484\,
            I => \N__5479\
        );

    \I__613\ : Span4Mux_h
    port map (
            O => \N__5479\,
            I => \N__5476\
        );

    \I__612\ : Odrv4
    port map (
            O => \N__5476\,
            I => \inst_midgetv_core.B_18\
        );

    \I__611\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5457\
        );

    \I__610\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5457\
        );

    \I__609\ : InMux
    port map (
            O => \N__5471\,
            I => \N__5457\
        );

    \I__608\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5457\
        );

    \I__607\ : InMux
    port map (
            O => \N__5469\,
            I => \N__5448\
        );

    \I__606\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5448\
        );

    \I__605\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5448\
        );

    \I__604\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5448\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__5457\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa13b\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5448\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa13b\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__5443\,
            I => \N__5435\
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__5442\,
            I => \N__5431\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__5441\,
            I => \N__5428\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__5440\,
            I => \N__5425\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__5439\,
            I => \N__5422\
        );

    \I__596\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5416\
        );

    \I__595\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5416\
        );

    \I__594\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5411\
        );

    \I__593\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5411\
        );

    \I__592\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5408\
        );

    \I__591\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5401\
        );

    \I__590\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5401\
        );

    \I__589\ : InMux
    port map (
            O => \N__5421\,
            I => \N__5401\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__5416\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa31\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__5411\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa31\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__5408\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa31\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__5401\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa31\
        );

    \I__584\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5388\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__5391\,
            I => \N__5385\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__5388\,
            I => \N__5382\
        );

    \I__581\ : InMux
    port map (
            O => \N__5385\,
            I => \N__5379\
        );

    \I__580\ : Span4Mux_h
    port map (
            O => \N__5382\,
            I => \N__5376\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__5379\,
            I => \N__5373\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__5376\,
            I => \N__5370\
        );

    \I__577\ : Span4Mux_h
    port map (
            O => \N__5373\,
            I => \N__5367\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__5370\,
            I => \inst_midgetv_core.B_19\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__5367\,
            I => \inst_midgetv_core.B_19\
        );

    \I__574\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5359\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__572\ : Span4Mux_h
    port map (
            O => \N__5356\,
            I => \N__5353\
        );

    \I__571\ : Span4Mux_h
    port map (
            O => \N__5353\,
            I => \N__5349\
        );

    \I__570\ : InMux
    port map (
            O => \N__5352\,
            I => \N__5346\
        );

    \I__569\ : Span4Mux_v
    port map (
            O => \N__5349\,
            I => \N__5343\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__5346\,
            I => \N__5340\
        );

    \I__567\ : Odrv4
    port map (
            O => \N__5343\,
            I => \inst_midgetv_core.B_20\
        );

    \I__566\ : Odrv4
    port map (
            O => \N__5340\,
            I => \inst_midgetv_core.B_20\
        );

    \I__565\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__5332\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm4a\
        );

    \I__563\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5326\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__5326\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm11b\
        );

    \I__561\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5320\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__5320\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm11a\
        );

    \I__559\ : InMux
    port map (
            O => \N__5317\,
            I => \N__5314\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__5314\,
            I => \N__5310\
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__5313\,
            I => \N__5307\
        );

    \I__556\ : Span4Mux_v
    port map (
            O => \N__5310\,
            I => \N__5304\
        );

    \I__555\ : InMux
    port map (
            O => \N__5307\,
            I => \N__5301\
        );

    \I__554\ : Sp12to4
    port map (
            O => \N__5304\,
            I => \N__5298\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__5301\,
            I => \N__5295\
        );

    \I__552\ : Odrv12
    port map (
            O => \N__5298\,
            I => \inst_midgetv_core.B_12\
        );

    \I__551\ : Odrv4
    port map (
            O => \N__5295\,
            I => \inst_midgetv_core.B_12\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__5290\,
            I => \N__5287\
        );

    \I__549\ : InMux
    port map (
            O => \N__5287\,
            I => \N__5284\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__5284\,
            I => \inst_midgetv_core.inst_ucodepc.n5608\
        );

    \I__547\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__5278\,
            I => \inst_midgetv_core.inst_ucodepc.n5609\
        );

    \I__545\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5271\
        );

    \I__544\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5268\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__5271\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_0\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__5268\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_0\
        );

    \I__541\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5260\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__5260\,
            I => \N__5257\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__5257\,
            I => \N__5254\
        );

    \I__538\ : Span4Mux_h
    port map (
            O => \N__5254\,
            I => \N__5251\
        );

    \I__537\ : Span4Mux_h
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__536\ : Odrv4
    port map (
            O => \N__5248\,
            I => \inst_midgetv_core.QQ_0\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__5245\,
            I => \N__5241\
        );

    \I__534\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5236\
        );

    \I__533\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5236\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__5236\,
            I => \N__5233\
        );

    \I__531\ : Span4Mux_h
    port map (
            O => \N__5233\,
            I => \N__5230\
        );

    \I__530\ : Span4Mux_h
    port map (
            O => \N__5230\,
            I => \N__5227\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__5227\,
            I => \inst_midgetv_core.s_cyclecnt_1\
        );

    \I__528\ : CascadeMux
    port map (
            O => \N__5224\,
            I => \N__5220\
        );

    \I__527\ : CascadeMux
    port map (
            O => \N__5223\,
            I => \N__5217\
        );

    \I__526\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5214\
        );

    \I__525\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5211\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__5214\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_1\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__5211\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_1\
        );

    \I__522\ : CascadeMux
    port map (
            O => \N__5206\,
            I => \N__5203\
        );

    \I__521\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5200\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__5200\,
            I => \N__5197\
        );

    \I__519\ : Span4Mux_h
    port map (
            O => \N__5197\,
            I => \N__5194\
        );

    \I__518\ : Odrv4
    port map (
            O => \N__5194\,
            I => \inst_midgetv_core.QQ_1\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__5191\,
            I => \N__5188\
        );

    \I__516\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5184\
        );

    \I__515\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5181\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__5184\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_5\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__5181\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_5\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__5176\,
            I => \N__5173\
        );

    \I__511\ : InMux
    port map (
            O => \N__5173\,
            I => \N__5170\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__5170\,
            I => \N__5167\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__508\ : Odrv4
    port map (
            O => \N__5164\,
            I => \inst_midgetv_core.QQ_5\
        );

    \I__507\ : InMux
    port map (
            O => \N__5161\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_28\
        );

    \I__506\ : InMux
    port map (
            O => \N__5158\,
            I => \bfn_13_21_0_\
        );

    \I__505\ : InMux
    port map (
            O => \N__5155\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_30\
        );

    \I__504\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5133\
        );

    \I__503\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5133\
        );

    \I__502\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5133\
        );

    \I__501\ : InMux
    port map (
            O => \N__5149\,
            I => \N__5133\
        );

    \I__500\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5130\
        );

    \I__499\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5121\
        );

    \I__498\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5121\
        );

    \I__497\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5121\
        );

    \I__496\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5121\
        );

    \I__495\ : InMux
    port map (
            O => \N__5143\,
            I => \N__5100\
        );

    \I__494\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5100\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__5133\,
            I => \N__5092\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__5130\,
            I => \N__5087\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__5121\,
            I => \N__5087\
        );

    \I__490\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5078\
        );

    \I__489\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5078\
        );

    \I__488\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5078\
        );

    \I__487\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5078\
        );

    \I__486\ : InMux
    port map (
            O => \N__5116\,
            I => \N__5069\
        );

    \I__485\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5069\
        );

    \I__484\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5069\
        );

    \I__483\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5069\
        );

    \I__482\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5060\
        );

    \I__481\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5060\
        );

    \I__480\ : InMux
    port map (
            O => \N__5110\,
            I => \N__5060\
        );

    \I__479\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5060\
        );

    \I__478\ : InMux
    port map (
            O => \N__5108\,
            I => \N__5051\
        );

    \I__477\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5051\
        );

    \I__476\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5051\
        );

    \I__475\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5051\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__5100\,
            I => \N__5048\
        );

    \I__473\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5043\
        );

    \I__472\ : InMux
    port map (
            O => \N__5098\,
            I => \N__5043\
        );

    \I__471\ : InMux
    port map (
            O => \N__5097\,
            I => \N__5036\
        );

    \I__470\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5036\
        );

    \I__469\ : InMux
    port map (
            O => \N__5095\,
            I => \N__5036\
        );

    \I__468\ : Span4Mux_v
    port map (
            O => \N__5092\,
            I => \N__5033\
        );

    \I__467\ : Span4Mux_v
    port map (
            O => \N__5087\,
            I => \N__5030\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__5078\,
            I => \N__5025\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__5069\,
            I => \N__5025\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N__5020\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__5051\,
            I => \N__5020\
        );

    \I__462\ : Span4Mux_h
    port map (
            O => \N__5048\,
            I => \N__5017\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__5043\,
            I => \N__5012\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__5036\,
            I => \N__5012\
        );

    \I__459\ : Span4Mux_h
    port map (
            O => \N__5033\,
            I => \N__5009\
        );

    \I__458\ : Span4Mux_h
    port map (
            O => \N__5030\,
            I => \N__5004\
        );

    \I__457\ : Span4Mux_h
    port map (
            O => \N__5025\,
            I => \N__5004\
        );

    \I__456\ : Span4Mux_h
    port map (
            O => \N__5020\,
            I => \N__5001\
        );

    \I__455\ : Span4Mux_h
    port map (
            O => \N__5017\,
            I => \N__4998\
        );

    \I__454\ : Span4Mux_h
    port map (
            O => \N__5012\,
            I => \N__4995\
        );

    \I__453\ : Span4Mux_v
    port map (
            O => \N__5009\,
            I => \N__4990\
        );

    \I__452\ : Span4Mux_v
    port map (
            O => \N__5004\,
            I => \N__4990\
        );

    \I__451\ : Span4Mux_h
    port map (
            O => \N__5001\,
            I => \N__4987\
        );

    \I__450\ : Span4Mux_v
    port map (
            O => \N__4998\,
            I => \N__4982\
        );

    \I__449\ : Span4Mux_h
    port map (
            O => \N__4995\,
            I => \N__4982\
        );

    \I__448\ : Span4Mux_v
    port map (
            O => \N__4990\,
            I => \N__4979\
        );

    \I__447\ : Span4Mux_v
    port map (
            O => \N__4987\,
            I => \N__4976\
        );

    \I__446\ : Span4Mux_v
    port map (
            O => \N__4982\,
            I => \N__4973\
        );

    \I__445\ : Odrv4
    port map (
            O => \N__4979\,
            I => \inst_midgetv_core.s_alu_2\
        );

    \I__444\ : Odrv4
    port map (
            O => \N__4976\,
            I => \inst_midgetv_core.s_alu_2\
        );

    \I__443\ : Odrv4
    port map (
            O => \N__4973\,
            I => \inst_midgetv_core.s_alu_2\
        );

    \I__442\ : InMux
    port map (
            O => \N__4966\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_31\
        );

    \I__441\ : InMux
    port map (
            O => \N__4963\,
            I => \inst_midgetv_core.alu_carryout\
        );

    \I__440\ : CascadeMux
    port map (
            O => \N__4960\,
            I => \N__4957\
        );

    \I__439\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4954\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4954\,
            I => \inst_midgetv_core.inst_condcode.n2\
        );

    \I__437\ : CascadeMux
    port map (
            O => \N__4951\,
            I => \N__4947\
        );

    \I__436\ : CascadeMux
    port map (
            O => \N__4950\,
            I => \N__4944\
        );

    \I__435\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4941\
        );

    \I__434\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4938\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__4941\,
            I => \inst_midgetv_core.alu_carryout_THRU_CO\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4938\,
            I => \inst_midgetv_core.alu_carryout_THRU_CO\
        );

    \I__431\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4930\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4930\,
            I => \inst_midgetv_core.inst_condcode.n6\
        );

    \I__429\ : InMux
    port map (
            O => \N__4927\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_19\
        );

    \I__428\ : InMux
    port map (
            O => \N__4924\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_20\
        );

    \I__427\ : InMux
    port map (
            O => \N__4921\,
            I => \bfn_13_20_0_\
        );

    \I__426\ : InMux
    port map (
            O => \N__4918\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_22\
        );

    \I__425\ : InMux
    port map (
            O => \N__4915\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_23\
        );

    \I__424\ : InMux
    port map (
            O => \N__4912\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_24\
        );

    \I__423\ : InMux
    port map (
            O => \N__4909\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_25\
        );

    \I__422\ : InMux
    port map (
            O => \N__4906\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_26\
        );

    \I__421\ : InMux
    port map (
            O => \N__4903\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_27\
        );

    \I__420\ : InMux
    port map (
            O => \N__4900\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_10\
        );

    \I__419\ : InMux
    port map (
            O => \N__4897\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_11\
        );

    \I__418\ : InMux
    port map (
            O => \N__4894\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_12\
        );

    \I__417\ : InMux
    port map (
            O => \N__4891\,
            I => \bfn_13_19_0_\
        );

    \I__416\ : InMux
    port map (
            O => \N__4888\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_14\
        );

    \I__415\ : InMux
    port map (
            O => \N__4885\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_15\
        );

    \I__414\ : InMux
    port map (
            O => \N__4882\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_16\
        );

    \I__413\ : InMux
    port map (
            O => \N__4879\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_17\
        );

    \I__412\ : InMux
    port map (
            O => \N__4876\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_18\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__4873\,
            I => \N__4870\
        );

    \I__410\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4867\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4867\,
            I => \N__4864\
        );

    \I__408\ : Odrv4
    port map (
            O => \N__4864\,
            I => \inst_midgetv_core.QQ_2\
        );

    \I__407\ : InMux
    port map (
            O => \N__4861\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_2\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__4858\,
            I => \N__4855\
        );

    \I__405\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4852\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4852\,
            I => \N__4849\
        );

    \I__403\ : Odrv4
    port map (
            O => \N__4849\,
            I => \inst_midgetv_core.QQ_3\
        );

    \I__402\ : InMux
    port map (
            O => \N__4846\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_3\
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__4843\,
            I => \N__4840\
        );

    \I__400\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4837\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__4837\,
            I => \N__4834\
        );

    \I__398\ : Odrv4
    port map (
            O => \N__4834\,
            I => \inst_midgetv_core.QQ_4\
        );

    \I__397\ : InMux
    port map (
            O => \N__4831\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_4\
        );

    \I__396\ : InMux
    port map (
            O => \N__4828\,
            I => \bfn_13_18_0_\
        );

    \I__395\ : CascadeMux
    port map (
            O => \N__4825\,
            I => \N__4822\
        );

    \I__394\ : InMux
    port map (
            O => \N__4822\,
            I => \N__4819\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__4819\,
            I => \N__4816\
        );

    \I__392\ : Odrv12
    port map (
            O => \N__4816\,
            I => \inst_midgetv_core.QQ_6\
        );

    \I__391\ : InMux
    port map (
            O => \N__4813\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_6\
        );

    \I__390\ : InMux
    port map (
            O => \N__4810\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_7\
        );

    \I__389\ : InMux
    port map (
            O => \N__4807\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_8\
        );

    \I__388\ : InMux
    port map (
            O => \N__4804\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_9\
        );

    \I__387\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4798\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__4798\,
            I => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa07h\
        );

    \I__385\ : InMux
    port map (
            O => \N__4795\,
            I => \inst_midgetv_core.alu_carryin\
        );

    \I__384\ : InMux
    port map (
            O => \N__4792\,
            I => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_1\
        );

    \I__383\ : InMux
    port map (
            O => \N__4789\,
            I => \bfn_13_15_0_\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__4786\,
            I => \N__4783\
        );

    \I__381\ : InMux
    port map (
            O => \N__4783\,
            I => \N__4779\
        );

    \I__380\ : InMux
    port map (
            O => \N__4782\,
            I => \N__4776\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4779\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_6\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__4776\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_6\
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__4771\,
            I => \N__4768\
        );

    \I__376\ : InMux
    port map (
            O => \N__4768\,
            I => \N__4764\
        );

    \I__375\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4761\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__4764\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_3\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__4761\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_3\
        );

    \I__372\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4752\
        );

    \I__371\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4749\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__4752\,
            I => \N__4746\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__4749\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_2\
        );

    \I__368\ : Odrv4
    port map (
            O => \N__4746\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_2\
        );

    \I__367\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4737\
        );

    \I__366\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4734\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__4737\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_4\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__4734\,
            I => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_4\
        );

    \I__363\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4726\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__4726\,
            I => \inst_midgetv_core.inst_ucodepc.n28\
        );

    \I__361\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4720\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__4720\,
            I => \inst_midgetv_core.inst_ucodepc.n5610\
        );

    \I__359\ : InMux
    port map (
            O => \N__4717\,
            I => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_0\
        );

    \I__358\ : InMux
    port map (
            O => \N__4714\,
            I => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_1\
        );

    \I__357\ : InMux
    port map (
            O => \N__4711\,
            I => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_2\
        );

    \I__356\ : InMux
    port map (
            O => \N__4708\,
            I => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_3\
        );

    \I__355\ : InMux
    port map (
            O => \N__4705\,
            I => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_4\
        );

    \I__354\ : InMux
    port map (
            O => \N__4702\,
            I => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_5\
        );

    \I__353\ : InMux
    port map (
            O => \N__4699\,
            I => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_6\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__4696\,
            I => \N__4693\
        );

    \I__351\ : CascadeBuf
    port map (
            O => \N__4693\,
            I => \N__4690\
        );

    \I__350\ : CascadeMux
    port map (
            O => \N__4690\,
            I => \N__4687\
        );

    \I__349\ : CascadeBuf
    port map (
            O => \N__4687\,
            I => \N__4684\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__4684\,
            I => \N__4681\
        );

    \I__347\ : CascadeBuf
    port map (
            O => \N__4681\,
            I => \N__4678\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__4678\,
            I => \N__4675\
        );

    \I__345\ : CascadeBuf
    port map (
            O => \N__4675\,
            I => \N__4672\
        );

    \I__344\ : CascadeMux
    port map (
            O => \N__4672\,
            I => \N__4669\
        );

    \I__343\ : CascadeBuf
    port map (
            O => \N__4669\,
            I => \N__4666\
        );

    \I__342\ : CascadeMux
    port map (
            O => \N__4666\,
            I => \N__4663\
        );

    \I__341\ : CascadeBuf
    port map (
            O => \N__4663\,
            I => \N__4660\
        );

    \I__340\ : CascadeMux
    port map (
            O => \N__4660\,
            I => \N__4657\
        );

    \I__339\ : CascadeBuf
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__4654\,
            I => \N__4651\
        );

    \I__337\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4648\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__4648\,
            I => \N__4645\
        );

    \I__335\ : Span4Mux_s3_v
    port map (
            O => \N__4645\,
            I => \N__4642\
        );

    \I__334\ : Span4Mux_v
    port map (
            O => \N__4642\,
            I => \N__4639\
        );

    \I__333\ : Sp12to4
    port map (
            O => \N__4639\,
            I => \N__4636\
        );

    \I__332\ : Span12Mux_h
    port map (
            O => \N__4636\,
            I => \N__4633\
        );

    \I__331\ : Odrv12
    port map (
            O => \N__4633\,
            I => \inst_midgetv_core.Wai_8\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy8\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy16\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy24\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy32\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_7\,
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_5_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_13\,
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_21\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_29\,
            carryinitout => \bfn_13_21_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_genblk1_L_93_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__13357\,
            in1 => \N__13441\,
            in2 => \_gnd_net_\,
            in3 => \N__6973\,
            lcout => \inst_midgetv_core.Wai_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i3947_4_lut_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__11853\,
            in1 => \N__8236\,
            in2 => \N__11830\,
            in3 => \N__12751\,
            lcout => \inst_midgetv_core.inst_ucodepc.n5610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i35_3_lut_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8908\,
            in1 => \N__9757\,
            in2 => \_gnd_net_\,
            in3 => \N__12473\,
            lcout => \inst_midgetv_core.inst_ucodepc.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i3962_4_lut_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__4729\,
            in1 => \N__11418\,
            in2 => \N__11875\,
            in3 => \N__4723\,
            lcout => \inst_midgetv_core.inst_ucodepc.n5608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_r_rcntlsb_0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__11189\,
            in1 => \N__5275\,
            in2 => \_gnd_net_\,
            in3 => \N__12991\,
            lcout => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_0\,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_0\,
            clk => \N__13806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_r_rcntlsb_1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__12992\,
            in1 => \N__11179\,
            in2 => \N__5224\,
            in3 => \N__4717\,
            lcout => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_1\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_0\,
            carryout => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_1\,
            clk => \N__13806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_r_rcntlsb_2_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__12996\,
            in1 => \N__4755\,
            in2 => \N__11197\,
            in3 => \N__4714\,
            lcout => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_2\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_1\,
            carryout => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_2\,
            clk => \N__13806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_r_rcntlsb_3_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__12993\,
            in1 => \N__11183\,
            in2 => \N__4771\,
            in3 => \N__4711\,
            lcout => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_3\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_2\,
            carryout => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_3\,
            clk => \N__13806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_r_rcntlsb_4_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__12997\,
            in1 => \N__4741\,
            in2 => \N__11198\,
            in3 => \N__4708\,
            lcout => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_4\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_3\,
            carryout => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_4\,
            clk => \N__13806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_r_rcntlsb_5_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__12994\,
            in1 => \N__11187\,
            in2 => \N__5191\,
            in3 => \N__4705\,
            lcout => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_5\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_4\,
            carryout => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_5\,
            clk => \N__13806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_r_buserror_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13549\,
            in1 => \N__12990\,
            in2 => \_gnd_net_\,
            in3 => \N__4702\,
            lcout => \inst_midgetv_core.buserror\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_5\,
            carryout => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_6\,
            clk => \N__13806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_r_rcntlsb_6_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__12995\,
            in1 => \N__11188\,
            in2 => \N__4786\,
            in3 => \N__4699\,
            lcout => \inst_midgetv_core.inst_cyclecnt.dbg_rccnt_6\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_6\,
            carryout => \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_ccntcy_7\,
            clk => \N__13806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_r_rcrun_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10625\,
            in2 => \_gnd_net_\,
            in3 => \N__4789\,
            lcout => corerunning,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_c_qq_62_4.l_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4782\,
            in1 => \N__11168\,
            in2 => \_gnd_net_\,
            in3 => \N__10230\,
            lcout => \inst_midgetv_core.QQ_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_c_qq_62_1.l_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11166\,
            in1 => \N__4767\,
            in2 => \_gnd_net_\,
            in3 => \N__11770\,
            lcout => \inst_midgetv_core.QQ_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_c_qq_62_0.l_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4756\,
            in1 => \N__11165\,
            in2 => \_gnd_net_\,
            in3 => \N__11510\,
            lcout => \inst_midgetv_core.QQ_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1796_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010100000"
        )
    port map (
            in0 => \N__10980\,
            in1 => \N__10899\,
            in2 => \N__10837\,
            in3 => \N__10270\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm4a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_l_sa09_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7768\,
            in2 => \_gnd_net_\,
            in3 => \N__11169\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_c_qq_62_2.l_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4740\,
            in1 => \N__11167\,
            in2 => \_gnd_net_\,
            in3 => \N__10449\,
            lcout => \inst_midgetv_core.QQ_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1605_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101011"
        )
    port map (
            in0 => \N__8867\,
            in1 => \N__10955\,
            in2 => \N__10836\,
            in3 => \N__10887\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_l_sa07_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4801\,
            in2 => \_gnd_net_\,
            in3 => \N__11190\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa07\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1804_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000000000"
        )
    port map (
            in0 => \N__10829\,
            in1 => \N__10960\,
            in2 => \N__14391\,
            in3 => \N__10889\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm11a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1598_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100101"
        )
    port map (
            in0 => \N__11268\,
            in1 => \N__11105\,
            in2 => \N__11323\,
            in3 => \N__8337\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa07h\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1603_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__10823\,
            in1 => \N__10954\,
            in2 => \_gnd_net_\,
            in3 => \N__10886\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1606_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000011"
        )
    port map (
            in0 => \N__10888\,
            in1 => \N__10827\,
            in2 => \N__10981\,
            in3 => \N__8868\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa13b\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1604_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100010001"
        )
    port map (
            in0 => \N__10822\,
            in1 => \N__10953\,
            in2 => \_gnd_net_\,
            in3 => \N__10885\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1805_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010100000"
        )
    port map (
            in0 => \N__10956\,
            in1 => \N__10039\,
            in2 => \N__8872\,
            in3 => \N__10828\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm11b\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu_carryin.genblk1_genblk1_lb.l_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__8404\,
            in1 => \N__8253\,
            in2 => \N__7131\,
            in3 => \N__8756\,
            lcout => \inst_midgetv_core.sra_msb\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \inst_midgetv_core.inst_alu_carryin.genblk1_genblk1_prealucyin\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu_carryin.genblk1_genblk1_reglastshift_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12415\,
            in2 => \N__12136\,
            in3 => \N__12788\,
            lcout => \inst_midgetv_core.rlastshift\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu_carryin.genblk1_genblk1_prealucyin\,
            carryout => \inst_midgetv_core.alu_carryin\,
            clk => \N__13791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_0.l_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5095\,
            in1 => \N__5263\,
            in2 => \N__6565\,
            in3 => \N__4795\,
            lcout => \inst_midgetv_core.B_0\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.alu_carryin\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_1.l_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5098\,
            in1 => \N__6487\,
            in2 => \N__5206\,
            in3 => \N__4792\,
            lcout => \inst_midgetv_core.B_1\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_1\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_2.l_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5096\,
            in1 => \N__6874\,
            in2 => \N__4873\,
            in3 => \N__4861\,
            lcout => \inst_midgetv_core.B_2\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_2\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_3.l_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5099\,
            in1 => \N__6832\,
            in2 => \N__4858\,
            in3 => \N__4846\,
            lcout => \inst_midgetv_core.B_3\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_3\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_4.l_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5097\,
            in1 => \N__6802\,
            in2 => \N__4843\,
            in3 => \N__4831\,
            lcout => \inst_midgetv_core.B_4\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_4\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_4.y_THRU_CRY_0_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12906\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_5\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_5_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_5.l_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5105\,
            in1 => \N__6775\,
            in2 => \N__5176\,
            in3 => \N__4828\,
            lcout => \inst_midgetv_core.B_5\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_6.l_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5109\,
            in1 => \N__7081\,
            in2 => \N__4825\,
            in3 => \N__4813\,
            lcout => \inst_midgetv_core.B_6\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_6\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_7.l_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5106\,
            in1 => \N__10143\,
            in2 => \N__7486\,
            in3 => \N__4810\,
            lcout => \inst_midgetv_core.B_7\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_7\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_8.l_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5111\,
            in1 => \N__13266\,
            in2 => \N__7051\,
            in3 => \N__4807\,
            lcout => \inst_midgetv_core.B_8\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_8\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_9.l_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5107\,
            in1 => \N__6925\,
            in2 => \N__6892\,
            in3 => \N__4804\,
            lcout => \inst_midgetv_core.B_9\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_9\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_10.l_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5110\,
            in1 => \N__6969\,
            in2 => \N__7018\,
            in3 => \N__4900\,
            lcout => \inst_midgetv_core.B_10\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_10\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_11.l_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5108\,
            in1 => \N__6985\,
            in2 => \N__11736\,
            in3 => \N__4897\,
            lcout => \inst_midgetv_core.B_11\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_11\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_12.l_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5112\,
            in1 => \N__7264\,
            in2 => \N__7288\,
            in3 => \N__4894\,
            lcout => \inst_midgetv_core.B_12\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_12\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_13.l_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5113\,
            in1 => \N__8593\,
            in2 => \N__8620\,
            in3 => \N__4891\,
            lcout => \inst_midgetv_core.B_13\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_14.l_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5117\,
            in1 => \N__9571\,
            in2 => \N__9601\,
            in3 => \N__4888\,
            lcout => \inst_midgetv_core.B_14\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_14\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_15.l_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5114\,
            in1 => \N__9517\,
            in2 => \N__9547\,
            in3 => \N__4885\,
            lcout => \inst_midgetv_core.B_15\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_15\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_16.l_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5119\,
            in1 => \N__9323\,
            in2 => \N__8962\,
            in3 => \N__4882\,
            lcout => \inst_midgetv_core.B_16\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_16\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_17.l_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5115\,
            in1 => \N__7456\,
            in2 => \N__9508\,
            in3 => \N__4879\,
            lcout => \inst_midgetv_core.B_17\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_17\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_18.l_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5118\,
            in1 => \N__7429\,
            in2 => \N__7405\,
            in3 => \N__4876\,
            lcout => \inst_midgetv_core.B_18\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_18\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_19.l_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5116\,
            in1 => \N__7354\,
            in2 => \N__7381\,
            in3 => \N__4927\,
            lcout => \inst_midgetv_core.B_19\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_19\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_20.l_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5120\,
            in1 => \N__7726\,
            in2 => \N__7753\,
            in3 => \N__4924\,
            lcout => \inst_midgetv_core.B_20\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_20\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_21.l_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5144\,
            in1 => \N__7330\,
            in2 => \N__5962\,
            in3 => \N__4921\,
            lcout => \inst_midgetv_core.B_21\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_22.l_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5149\,
            in1 => \N__5911\,
            in2 => \N__5935\,
            in3 => \N__4918\,
            lcout => \inst_midgetv_core.B_22\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_22\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_23.l_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5145\,
            in1 => \N__6475\,
            in2 => \N__6451\,
            in3 => \N__4915\,
            lcout => \inst_midgetv_core.B_23\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_23\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_24.l_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5150\,
            in1 => \N__6421\,
            in2 => \N__6397\,
            in3 => \N__4912\,
            lcout => \inst_midgetv_core.B_24\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_24\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_25.l_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5146\,
            in1 => \N__7669\,
            in2 => \N__7696\,
            in3 => \N__4909\,
            lcout => \inst_midgetv_core.B_25\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_25\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_26.l_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5151\,
            in1 => \N__7639\,
            in2 => \N__7615\,
            in3 => \N__4906\,
            lcout => \inst_midgetv_core.B_26\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_26\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_27.l_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5147\,
            in1 => \N__7558\,
            in2 => \N__7585\,
            in3 => \N__4903\,
            lcout => \inst_midgetv_core.B_27\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_27\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_28.l_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5152\,
            in1 => \N__8095\,
            in2 => \N__8068\,
            in3 => \N__5161\,
            lcout => \inst_midgetv_core.B_28\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_28\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_29.l_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5143\,
            in1 => \N__7549\,
            in2 => \N__7231\,
            in3 => \N__5158\,
            lcout => \inst_midgetv_core.B_29\,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_30.l_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5148\,
            in1 => \N__7171\,
            in2 => \N__7195\,
            in3 => \N__5155\,
            lcout => \inst_midgetv_core.B_30\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_30\,
            carryout => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.b_31.l_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__5142\,
            in1 => \N__7100\,
            in2 => \N__7144\,
            in3 => \N__4966\,
            lcout => \inst_midgetv_core.B_31\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_alu.genblk1_inst.alucy_31\,
            carryout => \inst_midgetv_core.alu_carryout\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.alu_carryout_THRU_LUT4_0_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4963\,
            lcout => \inst_midgetv_core.alu_carryout_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_condcode.genblk1_tmp_raluF_31_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__4933\,
            in1 => \N__8676\,
            in2 => \N__4960\,
            in3 => \N__8568\,
            lcout => \inst_midgetv_core.raluF\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_condcode.INSTR_14__I_0_i2_3_lut_4_lut_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001110"
        )
    port map (
            in0 => \N__7142\,
            in1 => \N__7101\,
            in2 => \N__4951\,
            in3 => \N__8211\,
            lcout => \inst_midgetv_core.inst_condcode.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_condcode.INSTR_14__I_0_i6_3_lut_4_lut_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001110"
        )
    port map (
            in0 => \N__7102\,
            in1 => \N__7143\,
            in2 => \N__4950\,
            in3 => \N__8675\,
            lcout => \inst_midgetv_core.inst_condcode.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i3958_2_lut_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11267\,
            in2 => \_gnd_net_\,
            in3 => \N__7821\,
            lcout => \inst_midgetv_core.inst_ucodepc.n5609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i1_4_lut_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010111010"
        )
    port map (
            in0 => \N__11944\,
            in1 => \N__7882\,
            in2 => \N__5290\,
            in3 => \N__5281\,
            lcout => \inst_midgetv_core.mostofminx0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_genblk1_c_qq_10_0.l_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101111"
        )
    port map (
            in0 => \N__6580\,
            in1 => \N__5274\,
            in2 => \N__5245\,
            in3 => \N__11162\,
            lcout => \inst_midgetv_core.QQ_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.reg_d18_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7947\,
            in1 => \N__6261\,
            in2 => \N__6298\,
            in3 => \N__7989\,
            lcout => \inst_midgetv_core.s_cyclecnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13811\,
            ce => \N__9808\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_genblk1_c_qq_10_1.l_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011101"
        )
    port map (
            in0 => \N__5244\,
            in1 => \N__6504\,
            in2 => \N__5223\,
            in3 => \N__11163\,
            lcout => \inst_midgetv_core.QQ_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_cyclecnt.genblk1_genblk1_c_qq_62_3.l_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5187\,
            in1 => \N__11164\,
            in2 => \_gnd_net_\,
            in3 => \N__10356\,
            lcout => \inst_midgetv_core.QQ_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_0__r_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__10900\,
            in1 => \N__12465\,
            in2 => \N__10832\,
            in3 => \N__10006\,
            lcout => \inst_midgetv_core.ADR_O_0\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy1\,
            clk => \N__13807\,
            ce => \N__9735\,
            sr => \N__6678\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_1__r_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__11011\,
            in1 => \N__12750\,
            in2 => \N__10901\,
            in3 => \N__13169\,
            lcout => \inst_midgetv_core.ADR_O_1\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy1\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy2\,
            clk => \N__13807\,
            ce => \N__9735\,
            sr => \N__6678\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_2__r_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__9955\,
            in1 => \N__10880\,
            in2 => \N__14200\,
            in3 => \N__15198\,
            lcout => \ADR_O_2\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy2\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy3\,
            clk => \N__13807\,
            ce => \N__9735\,
            sr => \N__6678\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_3__r_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111110100000"
        )
    port map (
            in0 => \N__13058\,
            in1 => \N__14051\,
            in2 => \N__10902\,
            in3 => \N__10729\,
            lcout => \ADR_O_3\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy3\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy4\,
            clk => \N__13807\,
            ce => \N__9735\,
            sr => \N__6678\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_4__r_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__14476\,
            in1 => \N__10884\,
            in2 => \N__15131\,
            in3 => \N__5335\,
            lcout => \inst_midgetv_core.ADR_O_4\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy4\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy5\,
            clk => \N__13807\,
            ce => \N__9735\,
            sr => \N__6678\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_5__r_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__8764\,
            in1 => \N__15306\,
            in2 => \N__10982\,
            in3 => \N__6120\,
            lcout => \inst_midgetv_core.ADR_O_5\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy5\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy6\,
            clk => \N__13807\,
            ce => \N__9735\,
            sr => \N__6678\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_6__r_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__6121\,
            in1 => \N__10964\,
            in2 => \N__14291\,
            in3 => \N__8833\,
            lcout => \inst_midgetv_core.ADR_O_6\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy6\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy7\,
            clk => \N__13807\,
            ce => \N__9735\,
            sr => \N__6678\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_7__r_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__8467\,
            in1 => \N__13919\,
            in2 => \N__10983\,
            in3 => \N__6119\,
            lcout => \inst_midgetv_core.ADR_O_7\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy7\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy8\,
            clk => \N__13807\,
            ce => \N__9735\,
            sr => \N__6678\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_8__r_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__6056\,
            in1 => \N__14780\,
            in2 => \N__10984\,
            in3 => \N__8796\,
            lcout => \inst_midgetv_core.ADR_O_8\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy9\,
            clk => \N__13801\,
            ce => \N__9727\,
            sr => \N__6681\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_9__r_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__8440\,
            in1 => \N__14606\,
            in2 => \N__10986\,
            in3 => \N__6057\,
            lcout => \inst_midgetv_core.ADR_O_9\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy9\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy10\,
            clk => \N__13801\,
            ce => \N__9727\,
            sr => \N__6681\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_10__r_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__6055\,
            in1 => \N__14978\,
            in2 => \N__10985\,
            in3 => \N__8400\,
            lcout => \inst_midgetv_core.ADR_O_10\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy10\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy11\,
            clk => \N__13801\,
            ce => \N__9727\,
            sr => \N__6681\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_11__r_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110101010"
        )
    port map (
            in0 => \N__5329\,
            in1 => \N__14885\,
            in2 => \N__12989\,
            in3 => \N__5323\,
            lcout => \inst_midgetv_core.ADR_O_11\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy11\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy12\,
            clk => \N__13801\,
            ce => \N__9727\,
            sr => \N__6681\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_12__r_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__5466\,
            in1 => \N__5421\,
            in2 => \N__5313\,
            in3 => \N__8203\,
            lcout => \inst_midgetv_core.ADR_O_12\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy12\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy13\,
            clk => \N__13801\,
            ce => \N__9727\,
            sr => \N__6681\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_13__r_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__8677\,
            in1 => \N__5637\,
            in2 => \N__5439\,
            in3 => \N__5468\,
            lcout => \inst_midgetv_core.ADR_O_13\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy13\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy14\,
            clk => \N__13801\,
            ce => \N__9727\,
            sr => \N__6681\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_14__r_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__5467\,
            in1 => \N__5610\,
            in2 => \N__5441\,
            in3 => \N__8569\,
            lcout => \inst_midgetv_core.ADR_O_14\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy14\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy15\,
            clk => \N__13801\,
            ce => \N__9727\,
            sr => \N__6681\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_15__r_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__14334\,
            in1 => \N__5586\,
            in2 => \N__5440\,
            in3 => \N__5469\,
            lcout => \inst_midgetv_core.ADR_O_15\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy15\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy16\,
            clk => \N__13801\,
            ce => \N__9727\,
            sr => \N__6681\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_16__r_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__13141\,
            in1 => \N__5556\,
            in2 => \N__5442\,
            in3 => \N__5472\,
            lcout => \inst_midgetv_core.ADR_O_16\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy17\,
            clk => \N__13797\,
            ce => \N__9736\,
            sr => \N__6679\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_17__r_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__5470\,
            in1 => \N__5526\,
            in2 => \N__5443\,
            in3 => \N__15162\,
            lcout => \inst_midgetv_core.ADR_O_17\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy17\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy18\,
            clk => \N__13797\,
            ce => \N__9736\,
            sr => \N__6679\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_18__r_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__13104\,
            in1 => \N__5438\,
            in2 => \N__5503\,
            in3 => \N__5473\,
            lcout => \inst_midgetv_core.ADR_O_18\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy18\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy19\,
            clk => \N__13797\,
            ce => \N__9736\,
            sr => \N__6679\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_19__r_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__5471\,
            in1 => \N__5434\,
            in2 => \N__5391\,
            in3 => \N__14430\,
            lcout => \inst_midgetv_core.ADR_O_19\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy19\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy20\,
            clk => \N__13797\,
            ce => \N__9736\,
            sr => \N__6679\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_20__r_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__14386\,
            in1 => \N__5352\,
            in2 => \N__6061\,
            in3 => \N__6145\,
            lcout => \inst_midgetv_core.ADR_O_20\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy20\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy21\,
            clk => \N__13797\,
            ce => \N__9736\,
            sr => \N__6679\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_21__r_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__6143\,
            in1 => \N__5883\,
            in2 => \N__6063\,
            in3 => \N__13176\,
            lcout => \inst_midgetv_core.ADR_O_21\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy21\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy22\,
            clk => \N__13797\,
            ce => \N__9736\,
            sr => \N__6679\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_22__r_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__15197\,
            in1 => \N__5847\,
            in2 => \N__6062\,
            in3 => \N__6146\,
            lcout => \inst_midgetv_core.ADR_O_22\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy22\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy23\,
            clk => \N__13797\,
            ce => \N__9736\,
            sr => \N__6679\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_23__r_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__6144\,
            in1 => \N__5820\,
            in2 => \N__6064\,
            in3 => \N__13059\,
            lcout => \inst_midgetv_core.ADR_O_23\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy23\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy24\,
            clk => \N__13797\,
            ce => \N__9736\,
            sr => \N__6679\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_24__r_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__14465\,
            in1 => \N__6065\,
            in2 => \N__5796\,
            in3 => \N__6168\,
            lcout => \inst_midgetv_core.ADR_O_24\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy25\,
            clk => \N__13792\,
            ce => \N__9728\,
            sr => \N__6680\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_25__r_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__6165\,
            in1 => \N__5754\,
            in2 => \N__6088\,
            in3 => \N__8760\,
            lcout => \inst_midgetv_core.ADR_O_25\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy25\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy26\,
            clk => \N__13792\,
            ce => \N__9728\,
            sr => \N__6680\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_26__r_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__8829\,
            in1 => \N__5724\,
            in2 => \N__6091\,
            in3 => \N__6169\,
            lcout => \inst_midgetv_core.ADR_O_26\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy26\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy27\,
            clk => \N__13792\,
            ce => \N__9728\,
            sr => \N__6680\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_27__r_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__8465\,
            in1 => \N__6078\,
            in2 => \N__5694\,
            in3 => \N__6172\,
            lcout => \inst_midgetv_core.ADR_O_27\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy27\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy28\,
            clk => \N__13792\,
            ce => \N__9728\,
            sr => \N__6680\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_28__r_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__8797\,
            in1 => \N__5661\,
            in2 => \N__6092\,
            in3 => \N__6170\,
            lcout => \inst_midgetv_core.ADR_O_28\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy28\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy29\,
            clk => \N__13792\,
            ce => \N__9728\,
            sr => \N__6680\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_29__r_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__6166\,
            in1 => \N__6192\,
            in2 => \N__6089\,
            in3 => \N__8438\,
            lcout => \inst_midgetv_core.ADR_O_29\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy29\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy30\,
            clk => \N__13792\,
            ce => \N__9728\,
            sr => \N__6680\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_30__r_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__8416\,
            in1 => \N__8943\,
            in2 => \N__6093\,
            in3 => \N__6171\,
            lcout => \inst_midgetv_core.ADR_O_30\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy30\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy31\,
            clk => \N__13792\,
            ce => \N__9728\,
            sr => \N__6680\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_blk0_31__r_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__6167\,
            in1 => \N__11433\,
            in2 => \N__6090\,
            in3 => \N__8866\,
            lcout => \inst_midgetv_core.ADR_O_31\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy31\,
            carryout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_zcy32\,
            clk => \N__13792\,
            ce => \N__9728\,
            sr => \N__6680\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_rNE0_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5986\,
            lcout => \inst_midgetv_core.rzcy32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13789\,
            ce => \N__9726\,
            sr => \N__6682\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_21_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5930\,
            in2 => \N__5983\,
            in3 => \N__9460\,
            lcout => \inst_midgetv_core.INSTR_21\,
            ltout => \inst_midgetv_core.Di_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13786\,
            ce => \N__9918\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_21.l_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__7326\,
            in1 => \N__9301\,
            in2 => \N__5965\,
            in3 => \N__9124\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_22_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6470\,
            in2 => \N__5953\,
            in3 => \N__9461\,
            lcout => \inst_midgetv_core.INSTR_22\,
            ltout => \inst_midgetv_core.Di_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13786\,
            ce => \N__9918\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_22.l_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__5931\,
            in1 => \N__9302\,
            in2 => \N__5914\,
            in3 => \N__9125\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_23_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6419\,
            in2 => \N__5905\,
            in3 => \N__9462\,
            lcout => \inst_midgetv_core.INSTR_23\,
            ltout => \inst_midgetv_core.Di_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13786\,
            ce => \N__9918\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_23.l_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__6471\,
            in1 => \N__9303\,
            in2 => \N__6454\,
            in3 => \N__9126\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_24_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7691\,
            in2 => \N__6442\,
            in3 => \N__9463\,
            lcout => \inst_midgetv_core.INSTR_24\,
            ltout => \inst_midgetv_core.Di_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13786\,
            ce => \N__9918\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_24.l_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__6420\,
            in1 => \N__9304\,
            in2 => \N__6400\,
            in3 => \N__9127\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.genblk4_rWE_O_66_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__8935\,
            in1 => \N__11353\,
            in2 => \_gnd_net_\,
            in3 => \N__11417\,
            lcout => \WE_O\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13785\,
            ce => \N__6736\,
            sr => \N__6721\
        );

    \inst_midgetv_core.inst_wai.genblk1_L_2327_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__13344\,
            in1 => \N__13442\,
            in2 => \_gnd_net_\,
            in3 => \N__6924\,
            lcout => \inst_midgetv_core.Wai_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.leq0100.l_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7902\,
            in1 => \N__6216\,
            in2 => \N__8031\,
            in3 => \N__6312\,
            lcout => \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.instr0100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.rinx_7__I_0_i3_4_lut_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__7823\,
            in1 => \N__7877\,
            in2 => \N__6283\,
            in3 => \N__11322\,
            lcout => \inst_midgetv_core.minx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.rinx_7__I_0_i1_4_lut_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__7876\,
            in1 => \N__11107\,
            in2 => \N__6241\,
            in3 => \N__7822\,
            lcout => \inst_midgetv_core.minx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i1_4_lut_adj_51_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001100"
        )
    port map (
            in0 => \N__6586\,
            in1 => \N__10645\,
            in2 => \N__6517\,
            in3 => \N__8116\,
            lcout => \inst_midgetv_core.inst_ucodepc.illegal\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.i1_3_lut_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__6748\,
            in1 => \N__6708\,
            in2 => \_gnd_net_\,
            in3 => \N__11957\,
            lcout => \inst_midgetv_core.inst_progressctrl.n2764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.ctrlreg_we_I_7_2_lut_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__11956\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6696\,
            lcout => \inst_midgetv_core.inst_progressctrl.ctrlreg_we_N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.badalignment_I_0_70_4_lut_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001111"
        )
    port map (
            in0 => \N__11857\,
            in1 => \N__12492\,
            in2 => \N__10660\,
            in3 => \N__12727\,
            lcout => \inst_midgetv_core.inst_progressctrl.badalignment\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_cmb_sa14_or_nCORERUNNING_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6697\,
            in2 => \_gnd_net_\,
            in3 => \N__10646\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_nsa14_or_nCORERUNNING\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_0_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6617\,
            in2 => \N__6505\,
            in3 => \N__9375\,
            lcout => \inst_midgetv_core.INSTR_0\,
            ltout => \inst_midgetv_core.Di_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13812\,
            ce => \N__9876\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_0.l_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__6579\,
            in1 => \N__9247\,
            in2 => \N__6568\,
            in3 => \N__9013\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_1_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__6540\,
            in1 => \N__11508\,
            in2 => \_gnd_net_\,
            in3 => \N__9376\,
            lcout => \inst_midgetv_core.INSTR_1\,
            ltout => \inst_midgetv_core.Di_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13812\,
            ce => \N__9876\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_1.l_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000011100"
        )
    port map (
            in0 => \N__9197\,
            in1 => \N__9012\,
            in2 => \N__6508\,
            in3 => \N__6503\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_2_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__10557\,
            in1 => \_gnd_net_\,
            in2 => \N__11781\,
            in3 => \N__9377\,
            lcout => \inst_midgetv_core.INSTR_2\,
            ltout => \inst_midgetv_core.Di_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13812\,
            ce => \N__9876\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_2.l_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__11509\,
            in1 => \N__9248\,
            in2 => \N__6877\,
            in3 => \N__9015\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_3_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10447\,
            in2 => \N__6862\,
            in3 => \N__9378\,
            lcout => \inst_midgetv_core.INSTR_3\,
            ltout => \inst_midgetv_core.Di_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13812\,
            ce => \N__9876\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_3.l_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000011100"
        )
    port map (
            in0 => \N__9198\,
            in1 => \N__9014\,
            in2 => \N__6835\,
            in3 => \N__11769\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_4_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10354\,
            in2 => \N__6820\,
            in3 => \N__9379\,
            lcout => \inst_midgetv_core.INSTR_4\,
            ltout => \inst_midgetv_core.Di_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13808\,
            ce => \N__9901\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_4.l_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000011010"
        )
    port map (
            in0 => \N__9081\,
            in1 => \N__9254\,
            in2 => \N__6805\,
            in3 => \N__10448\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_5_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__6790\,
            in1 => \N__10228\,
            in2 => \_gnd_net_\,
            in3 => \N__9380\,
            lcout => \inst_midgetv_core.INSTR_5\,
            ltout => \inst_midgetv_core.Di_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13808\,
            ce => \N__9901\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_5.l_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011010010"
        )
    port map (
            in0 => \N__9082\,
            in1 => \N__10355\,
            in2 => \N__6778\,
            in3 => \N__9255\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_6_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10132\,
            in2 => \N__6763\,
            in3 => \N__9381\,
            lcout => \inst_midgetv_core.INSTR_6\,
            ltout => \inst_midgetv_core.Di_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13808\,
            ce => \N__9901\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_6.l_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010110100"
        )
    port map (
            in0 => \N__10229\,
            in1 => \N__9109\,
            in2 => \N__7084\,
            in3 => \N__9256\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_8_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__9445\,
            in1 => \N__6913\,
            in2 => \N__8887\,
            in3 => \N__7069\,
            lcout => \inst_midgetv_core.INSTR_8\,
            ltout => \inst_midgetv_core.Di_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13808\,
            ce => \N__9901\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_8.l_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011010010"
        )
    port map (
            in0 => \N__9083\,
            in1 => \N__13258\,
            in2 => \N__7054\,
            in3 => \N__9257\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_10_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11722\,
            in2 => \N__7036\,
            in3 => \N__9419\,
            lcout => \inst_midgetv_core.INSTR_10\,
            ltout => \inst_midgetv_core.Di_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13802\,
            ce => \N__9899\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_10.l_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__6962\,
            in1 => \N__9262\,
            in2 => \N__7021\,
            in3 => \N__9087\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_11_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7280\,
            in2 => \N__7003\,
            in3 => \N__9420\,
            lcout => \inst_midgetv_core.INSTR_11\,
            ltout => \inst_midgetv_core.Di_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13802\,
            ce => \N__9899\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_11.l_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__11723\,
            in1 => \N__9263\,
            in2 => \N__6988\,
            in3 => \N__9088\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_9_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6961\,
            in2 => \N__6943\,
            in3 => \N__9418\,
            lcout => \inst_midgetv_core.INSTR_9\,
            ltout => \inst_midgetv_core.Di_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13802\,
            ce => \N__9899\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_9.l_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000011100"
        )
    port map (
            in0 => \N__9249\,
            in1 => \N__9086\,
            in2 => \N__6928\,
            in3 => \N__6914\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_12_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8606\,
            in2 => \N__7306\,
            in3 => \N__9421\,
            lcout => \inst_midgetv_core.INSTR_12\,
            ltout => \inst_midgetv_core.Di_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13802\,
            ce => \N__9899\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_12.l_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__7281\,
            in1 => \N__9264\,
            in2 => \N__7267\,
            in3 => \N__9089\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_29_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7187\,
            in2 => \N__7252\,
            in3 => \N__9423\,
            lcout => \inst_midgetv_core.FUNC7_4\,
            ltout => \inst_midgetv_core.Di_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13798\,
            ce => \N__9911\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_29.l_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000011010"
        )
    port map (
            in0 => \N__9085\,
            in1 => \N__9259\,
            in2 => \N__7234\,
            in3 => \N__7544\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_30_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7126\,
            in2 => \N__7216\,
            in3 => \N__9424\,
            lcout => \inst_midgetv_core.FUNC7_5\,
            ltout => \inst_midgetv_core.Di_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13798\,
            ce => \N__9911\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_30.l_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__7188\,
            in1 => \N__9260\,
            in2 => \N__7174\,
            in3 => \N__9118\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_31_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__11641\,
            in1 => \N__7159\,
            in2 => \_gnd_net_\,
            in3 => \N__9425\,
            lcout => \inst_midgetv_core.FUNC7_6\,
            ltout => \inst_midgetv_core.Di_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13798\,
            ce => \N__9911\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_31.l_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__7127\,
            in1 => \N__9261\,
            in2 => \N__7105\,
            in3 => \N__9119\,
            lcout => \inst_midgetv_core.A31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_7_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__7504\,
            in1 => \N__13265\,
            in2 => \_gnd_net_\,
            in3 => \N__9422\,
            lcout => \inst_midgetv_core.INSTR_7\,
            ltout => \inst_midgetv_core.Di_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13798\,
            ce => \N__9911\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_7.l_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000011010"
        )
    port map (
            in0 => \N__9084\,
            in1 => \N__9258\,
            in2 => \N__7489\,
            in3 => \N__10142\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_17_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__9430\,
            in1 => \N__7474\,
            in2 => \_gnd_net_\,
            in3 => \N__7427\,
            lcout => \inst_midgetv_core.INSTR_17\,
            ltout => \inst_midgetv_core.Di_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13793\,
            ce => \N__9898\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_17.l_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000011100"
        )
    port map (
            in0 => \N__9253\,
            in1 => \N__9114\,
            in2 => \N__7459\,
            in3 => \N__9507\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_18_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__9431\,
            in1 => \N__7444\,
            in2 => \_gnd_net_\,
            in3 => \N__7376\,
            lcout => \inst_midgetv_core.INSTR_18\,
            ltout => \inst_midgetv_core.Di_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13793\,
            ce => \N__9898\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_18.l_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__7428\,
            in1 => \N__9294\,
            in2 => \N__7408\,
            in3 => \N__9115\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_19_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100100"
        )
    port map (
            in0 => \N__7393\,
            in1 => \N__7748\,
            in2 => \N__9455\,
            in3 => \_gnd_net_\,
            lcout => \inst_midgetv_core.INSTR_19\,
            ltout => \inst_midgetv_core.Di_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13793\,
            ce => \N__9898\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_19.l_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__7377\,
            in1 => \N__9295\,
            in2 => \N__7357\,
            in3 => \N__9116\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_20_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__9435\,
            in1 => \N__7345\,
            in2 => \_gnd_net_\,
            in3 => \N__7325\,
            lcout => \inst_midgetv_core.INSTR_20\,
            ltout => \inst_midgetv_core.Di_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13793\,
            ce => \N__9898\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_20.l_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__7749\,
            in1 => \N__9296\,
            in2 => \N__7729\,
            in3 => \N__9117\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_25_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7637\,
            in2 => \N__7717\,
            in3 => \N__9456\,
            lcout => \inst_midgetv_core.FUNC7_0\,
            ltout => \inst_midgetv_core.Di_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13790\,
            ce => \N__9919\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_25.l_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000011010"
        )
    port map (
            in0 => \N__9120\,
            in1 => \N__9297\,
            in2 => \N__7699\,
            in3 => \N__7695\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_26_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7580\,
            in2 => \N__7657\,
            in3 => \N__9457\,
            lcout => \inst_midgetv_core.FUNC7_1\,
            ltout => \inst_midgetv_core.Di_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13790\,
            ce => \N__9919\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_26.l_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__7638\,
            in1 => \N__9298\,
            in2 => \N__7618\,
            in3 => \N__9122\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_27_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8090\,
            in2 => \N__7603\,
            in3 => \N__9458\,
            lcout => \inst_midgetv_core.FUNC7_2\,
            ltout => \inst_midgetv_core.Di_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13790\,
            ce => \N__9919\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_27.l_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__7581\,
            in1 => \N__9299\,
            in2 => \N__7561\,
            in3 => \N__9123\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_28_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7545\,
            in2 => \N__7525\,
            in3 => \N__9459\,
            lcout => \inst_midgetv_core.FUNC7_3\,
            ltout => \inst_midgetv_core.Di_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13790\,
            ce => \N__9919\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_28.l_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__8091\,
            in1 => \N__9300\,
            in2 => \N__8071\,
            in3 => \N__9121\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.rinx_1__I_0_4_lut_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__7825\,
            in1 => \N__7869\,
            in2 => \N__8053\,
            in3 => \N__8149\,
            lcout => \inst_midgetv_core.minx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.rinx_7__I_0_i4_4_lut_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__7873\,
            in1 => \N__8212\,
            in2 => \N__8011\,
            in3 => \N__7826\,
            lcout => \inst_midgetv_core.minx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.usedinx_or_RST_I_notcorerunning_I_0_2_lut_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10650\,
            in2 => \_gnd_net_\,
            in3 => \N__11202\,
            lcout => \inst_midgetv_core.inst_ucodepc.usedinx_or_RST_I_notcorerunning\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.rinx_7__I_0_i6_4_lut_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__7874\,
            in1 => \N__7774\,
            in2 => \N__7966\,
            in3 => \N__7827\,
            lcout => \inst_midgetv_core.minx_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.rinx_7__I_0_i2_4_lut_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__8341\,
            in1 => \N__7921\,
            in2 => \N__7881\,
            in3 => \N__7824\,
            lcout => \inst_midgetv_core.minx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.rinx_7__I_0_i5_4_lut_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__7875\,
            in1 => \N__8131\,
            in2 => \N__7843\,
            in3 => \N__7828\,
            lcout => \inst_midgetv_core.minx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i1_3_lut_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__11256\,
            in1 => \N__8143\,
            in2 => \_gnd_net_\,
            in3 => \N__8561\,
            lcout => \inst_midgetv_core.inst_ucodepc.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_l_sa09h_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100011001"
        )
    port map (
            in0 => \N__11319\,
            in1 => \N__11252\,
            in2 => \N__8515\,
            in3 => \N__11108\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa09h\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i3950_4_lut_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__11110\,
            in1 => \N__8137\,
            in2 => \N__11266\,
            in3 => \N__8340\,
            lcout => \inst_midgetv_core.inst_ucodepc.n5603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i29_3_lut_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__8339\,
            in1 => \N__8511\,
            in2 => \_gnd_net_\,
            in3 => \N__11109\,
            lcout => \inst_midgetv_core.inst_ucodepc.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i255_4_lut_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__8510\,
            in1 => \N__11320\,
            in2 => \N__8415\,
            in3 => \N__8338\,
            lcout => \inst_midgetv_core.inst_ucodepc.dinx_1_N_145_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i3956_4_lut_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__11084\,
            in1 => \N__11245\,
            in2 => \N__8514\,
            in3 => \N__8666\,
            lcout => \inst_midgetv_core.inst_ucodepc.n5613\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i1545_4_lut_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__11083\,
            in1 => \N__11244\,
            in2 => \N__8513\,
            in3 => \N__8322\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk2_illegal_a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i2_4_lut_adj_50_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__8122\,
            in1 => \N__11300\,
            in2 => \N__8110\,
            in3 => \N__8521\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i1_4_lut_adj_49_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101000"
        )
    port map (
            in0 => \N__8716\,
            in1 => \N__8101\,
            in2 => \N__8266\,
            in3 => \N__8347\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i2_4_lut_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__11082\,
            in1 => \N__11243\,
            in2 => \N__11315\,
            in3 => \N__8321\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk1_checkfunct7_N_286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i256_4_lut_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000011100"
        )
    port map (
            in0 => \N__8664\,
            in1 => \N__8559\,
            in2 => \N__8336\,
            in3 => \N__8190\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i3967_4_lut_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110011"
        )
    port map (
            in0 => \N__8194\,
            in1 => \N__8473\,
            in2 => \N__8281\,
            in3 => \N__8899\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n5605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i1_4_lut_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100000000"
        )
    port map (
            in0 => \N__11242\,
            in1 => \N__11085\,
            in2 => \N__8512\,
            in3 => \N__8320\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i1_2_lut_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11081\,
            in2 => \_gnd_net_\,
            in3 => \N__8663\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n2575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_mimux.genblk1_sa00mod_r_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9679\,
            in1 => \N__10666\,
            in2 => \_gnd_net_\,
            in3 => \N__13615\,
            lcout => \inst_midgetv_core.inst_mimux.genblk1_sa00mod\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i4_4_lut_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__8466\,
            in1 => \N__8439\,
            in2 => \N__8414\,
            in3 => \N__8353\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i3_4_lut_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8319\,
            in1 => \N__11241\,
            in2 => \N__8204\,
            in3 => \N__8277\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk1_checkfunct7_N_281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_condcode.INSTR_14__I_0_32_i7_4_lut_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__8196\,
            in1 => \N__8257\,
            in2 => \N__8158\,
            in3 => \N__8560\,
            lcout => \inst_midgetv_core.is_brcond\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \STB_O_I_0_2_lut_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11795\,
            in2 => \_gnd_net_\,
            in3 => \N__13545\,
            lcout => \uart_ACK_O\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_condcode.i3953_3_lut_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__8224\,
            in1 => \N__8195\,
            in2 => \_gnd_net_\,
            in3 => \N__8665\,
            lcout => \inst_midgetv_core.inst_condcode.n5618\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i9_4_lut_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13130\,
            in1 => \N__10019\,
            in2 => \N__8701\,
            in3 => \N__8707\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.genblk1_illegal_rs1_rd_N_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_inputmux.genblk1_ireg__i1_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__10662\,
            in1 => \N__8893\,
            in2 => \N__10593\,
            in3 => \N__8886\,
            lcout => \rDee_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i5_4_lut_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__8849\,
            in1 => \N__8825\,
            in2 => \N__8795\,
            in3 => \N__8749\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i7_4_lut_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10742\,
            in1 => \N__14324\,
            in2 => \N__10262\,
            in3 => \N__15146\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.inst_illegalop.i6_4_lut_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9980\,
            in1 => \N__13094\,
            in2 => \N__14420\,
            in3 => \N__11033\,
            lcout => \inst_midgetv_core.inst_ucodepc.inst_illegalop.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_13_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9599\,
            in2 => \N__8692\,
            in3 => \N__9426\,
            lcout => \inst_midgetv_core.INSTR_13\,
            ltout => \inst_midgetv_core.Di_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13799\,
            ce => \N__9900\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_13.l_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000011100"
        )
    port map (
            in0 => \N__9293\,
            in1 => \N__9110\,
            in2 => \N__8623\,
            in3 => \N__8619\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_14_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9542\,
            in2 => \N__8584\,
            in3 => \N__9427\,
            lcout => \inst_midgetv_core.INSTR_14\,
            ltout => \inst_midgetv_core.Di_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13799\,
            ce => \N__9900\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_14.l_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__9600\,
            in1 => \N__9250\,
            in2 => \N__9574\,
            in3 => \N__9111\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC15_0_15_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9324\,
            in2 => \N__9562\,
            in3 => \N__9428\,
            lcout => \inst_midgetv_core.INSTR_15\,
            ltout => \inst_midgetv_core.Di_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13799\,
            ce => \N__9900\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_15.l_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__9543\,
            in1 => \N__9251\,
            in2 => \N__9520\,
            in3 => \N__9112\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_opreg.genblk1_OpC31_16_16_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9506\,
            in2 => \N__9481\,
            in3 => \N__9429\,
            lcout => \inst_midgetv_core.INSTR_16\,
            ltout => \inst_midgetv_core.Di_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13799\,
            ce => \N__9900\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_alu.genblk1_inst.a_16.l_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100110000"
        )
    port map (
            in0 => \N__9325\,
            in1 => \N__9252\,
            in2 => \N__9130\,
            in3 => \N__9113\,
            lcout => \inst_midgetv_core.inst_alu.genblk1_inst.A_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.i1_2_lut_3_lut_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__11373\,
            in1 => \N__8939\,
            in2 => \_gnd_net_\,
            in3 => \N__11345\,
            lcout => \inst_midgetv_core.inst_progressctrl.n4_adj_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d31_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__12325\,
            in1 => \N__12262\,
            in2 => \N__12399\,
            in3 => \N__12202\,
            lcout => \inst_midgetv_core.sa29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d15_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__12204\,
            in1 => \N__12327\,
            in2 => \N__12273\,
            in3 => \N__12392\,
            lcout => \inst_midgetv_core.is_valid_instrhigh\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.progress_ucode_I_0_4_lut_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011100"
        )
    port map (
            in0 => \N__13538\,
            in1 => \N__11964\,
            in2 => \N__10711\,
            in3 => \N__9742\,
            lcout => \inst_midgetv_core.progress_ucode\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d34_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__12203\,
            in1 => \N__12326\,
            in2 => \N__12272\,
            in3 => \N__12391\,
            lcout => \inst_midgetv_core.sa33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.i3968_4_lut_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11823\,
            in1 => \N__11846\,
            in2 => \N__9772\,
            in3 => \N__11868\,
            lcout => \inst_midgetv_core.inst_ucodepc.n5624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.i1_2_lut_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__9748\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12789\,
            lcout => \inst_midgetv_core.inst_progressctrl.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.blka_l_en_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10686\,
            lcout => \inst_midgetv_core.inst_progressctrl.blka_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.i1_4_lut_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__13537\,
            in1 => \N__11905\,
            in2 => \N__12793\,
            in3 => \N__11887\,
            lcout => \inst_midgetv_core.enaQ\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d08_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100100000"
        )
    port map (
            in0 => \N__12274\,
            in1 => \N__12208\,
            in2 => \N__12334\,
            in3 => \N__12400\,
            lcout => \inst_midgetv_core.sa00\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_L_2319_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__13330\,
            in1 => \N__10037\,
            in2 => \N__13430\,
            in3 => \N__10045\,
            lcout => \inst_midgetv_core.Wai_0\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \inst_midgetv_core.inst_wai.genblk1_waicy0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_L_2321_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__11743\,
            in1 => \N__13413\,
            in2 => \N__11041\,
            in3 => \N__13332\,
            lcout => \inst_midgetv_core.Wai_1\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_wai.genblk1_waicy0\,
            carryout => \inst_midgetv_core.inst_wai.genblk1_waicy1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_L_2322_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__13331\,
            in1 => \N__9987\,
            in2 => \N__13431\,
            in3 => \N__10453\,
            lcout => \inst_midgetv_core.Wai_2\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_wai.genblk1_waicy1\,
            carryout => \inst_midgetv_core.inst_wai.genblk1_waicy2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_L_2323_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__10360\,
            in1 => \N__13417\,
            in2 => \N__10762\,
            in3 => \N__13329\,
            lcout => \inst_midgetv_core.Wai_3\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_wai.genblk1_waicy2\,
            carryout => \inst_midgetv_core.inst_wai.genblk1_waicy3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_L_2324_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__13328\,
            in1 => \N__10269\,
            in2 => \N__13432\,
            in3 => \N__10240\,
            lcout => \inst_midgetv_core.Wai_4\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_wai.genblk1_waicy3\,
            carryout => \inst_midgetv_core.inst_wai.genblk1_waicy4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_L_2325_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011111110"
        )
    port map (
            in0 => \N__10144\,
            in1 => \N__13421\,
            in2 => \N__13365\,
            in3 => \N__10111\,
            lcout => \inst_midgetv_core.Wai_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_L_2318_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13327\,
            in1 => \N__12115\,
            in2 => \_gnd_net_\,
            in3 => \N__11534\,
            lcout => \inst_midgetv_core.inst_wai.genblk1_preWai0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1788_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__10996\,
            in1 => \N__10904\,
            in2 => \N__14390\,
            in3 => \N__10038\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm0a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1792_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001000000"
        )
    port map (
            in0 => \N__10903\,
            in1 => \N__10997\,
            in2 => \N__9991\,
            in3 => \N__10815\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm2a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.we_I_0_2_lut_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__12576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10717\,
            lcout => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrb.we\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1599_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100101111"
        )
    port map (
            in0 => \N__11321\,
            in1 => \N__11269\,
            in2 => \N__11203\,
            in3 => \N__11106\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_sa08\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1790_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010100000"
        )
    port map (
            in0 => \N__10998\,
            in1 => \N__10905\,
            in2 => \N__10831\,
            in3 => \N__11037\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm1a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_immexp_zfind_q.genblk1_L_1794_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010100000"
        )
    port map (
            in0 => \N__10999\,
            in1 => \N__10906\,
            in2 => \N__10830\,
            in3 => \N__10758\,
            lcout => \inst_midgetv_core.inst_immexp_zfind_q.genblk1_imm3a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.blka_r_bsel0_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000011100000100"
        )
    port map (
            in0 => \N__12117\,
            in1 => \N__12479\,
            in2 => \N__12070\,
            in3 => \N__12731\,
            lcout => \inst_midgetv_core.bmask_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13814\,
            ce => \N__12028\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.genblk6_l_iwe_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11560\,
            in1 => \N__10704\,
            in2 => \N__10687\,
            in3 => \N__10661\,
            lcout => \inst_midgetv_core.iwe\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.blka_r_bsel3_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000100000111"
        )
    port map (
            in0 => \N__12116\,
            in1 => \N__12478\,
            in2 => \N__12069\,
            in3 => \N__12730\,
            lcout => \inst_midgetv_core.bmask_3\,
            ltout => \inst_midgetv_core.inst_progressctrl.blka_cmb_bsel_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13814\,
            ce => \N__12028\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.blka_r_asel3_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10597\,
            in3 => \_gnd_net_\,
            lcout => \SEL_O_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13814\,
            ce => \N__12028\,
            sr => \_gnd_net_\
        );

    \i_LEDs.LED3_26_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__10594\,
            in1 => \N__11610\,
            in2 => \_gnd_net_\,
            in3 => \N__10561\,
            lcout => \LED3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13810\,
            ce => \N__11593\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_genblk1_genblk1_L_95_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__13361\,
            in1 => \N__13449\,
            in2 => \_gnd_net_\,
            in3 => \N__11737\,
            lcout => \inst_midgetv_core.Wai_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i_LEDs.bluesource_is_uart_25_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__11471\,
            in1 => \N__11650\,
            in2 => \N__11611\,
            in3 => \N__11637\,
            lcout => bluesource_is_uart,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i_LEDs.i1_2_lut_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11606\,
            in2 => \_gnd_net_\,
            in3 => \N__11470\,
            lcout => \i_LEDs.n2766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1538_2_lut_3_lut_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__13534\,
            in1 => \N__11794\,
            in2 => \_gnd_net_\,
            in3 => \N__11528\,
            lcout => \ACK_I\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_ACK_O_I_0_2_lut_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11802\,
            in2 => \_gnd_net_\,
            in3 => \N__11536\,
            lcout => n2345,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i_BBUART.STB_I_I_0_2_lut_3_lut_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11559\,
            in1 => \N__13521\,
            in2 => \_gnd_net_\,
            in3 => \N__11803\,
            lcout => \i_BBUART.usartTX_N_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i_LEDs.i2_3_lut_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11558\,
            in1 => \N__13520\,
            in2 => \_gnd_net_\,
            in3 => \N__11535\,
            lcout => \LED1_N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.genblk3_rSTB_O_64_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__11449\,
            in1 => \N__13533\,
            in2 => \N__11443\,
            in3 => \N__11426\,
            lcout => \STB_O\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13794\,
            ce => 'H',
            sr => \N__11971\
        );

    \inst_midgetv_core.inst_progressctrl.genblk3_rsram_stb_65_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__11425\,
            in1 => \N__13565\,
            in2 => \N__11380\,
            in3 => \N__11352\,
            lcout => \inst_midgetv_core.sram_stb\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13794\,
            ce => 'H',
            sr => \N__11971\
        );

    \CONSTANT_ZERO_LUT4_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ZERO_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d33_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100010010000"
        )
    port map (
            in0 => \N__12248\,
            in1 => \N__12172\,
            in2 => \N__12389\,
            in3 => \N__12304\,
            lcout => \inst_midgetv_core.sa32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucodepc.sa32_I_0_2_lut_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11901\,
            in2 => \_gnd_net_\,
            in3 => \N__11886\,
            lcout => \inst_midgetv_core.inst_ucodepc.maybranch_N_253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d32_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__12305\,
            in1 => \N__12375\,
            in2 => \N__12198\,
            in3 => \N__12250\,
            lcout => \inst_midgetv_core.sa30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d14_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__12249\,
            in1 => \N__12176\,
            in2 => \N__12390\,
            in3 => \N__12306\,
            lcout => \inst_midgetv_core.sa37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d38_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__12307\,
            in1 => \N__12371\,
            in2 => \N__12199\,
            in3 => \N__12247\,
            lcout => \inst_midgetv_core.sa40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.blka_l_usedefault_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101101"
        )
    port map (
            in0 => \N__11812\,
            in1 => \N__13299\,
            in2 => \N__12111\,
            in3 => \N__13390\,
            lcout => \inst_midgetv_core.inst_progressctrl.blka_usedefault\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d35_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000010"
        )
    port map (
            in0 => \N__12369\,
            in1 => \N__12312\,
            in2 => \N__12200\,
            in3 => \N__12242\,
            lcout => \inst_midgetv_core.sa34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_L_2320_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13298\,
            in1 => \N__11811\,
            in2 => \_gnd_net_\,
            in3 => \N__11801\,
            lcout => \inst_midgetv_core.inst_wai.genblk1_preWai1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d09_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000010000"
        )
    port map (
            in0 => \N__12241\,
            in1 => \N__12180\,
            in2 => \N__12324\,
            in3 => \N__12368\,
            lcout => \inst_midgetv_core.s_alu_carryin_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d21_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000111111"
        )
    port map (
            in0 => \N__12370\,
            in1 => \N__12313\,
            in2 => \N__12201\,
            in3 => \N__12243\,
            lcout => \inst_midgetv_core.s_shift_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ucode.genblk1_inst_2ebr.cmb_d10_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100000"
        )
    port map (
            in0 => \N__12367\,
            in1 => \N__12311\,
            in2 => \N__12261\,
            in3 => \N__12197\,
            lcout => \inst_midgetv_core.s_alu_carryin_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.blka_r_bsel1_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000011100000001"
        )
    port map (
            in0 => \N__12102\,
            in1 => \N__12495\,
            in2 => \N__12058\,
            in3 => \N__12726\,
            lcout => \inst_midgetv_core.bmask_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13822\,
            ce => \N__12027\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_progressctrl.blka_r_bsel2_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000010000000111"
        )
    port map (
            in0 => \N__12118\,
            in1 => \N__12494\,
            in2 => \N__12068\,
            in3 => \N__12725\,
            lcout => \inst_midgetv_core.bmask_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13819\,
            ce => \N__12026\,
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_shiftcounter.genblk1_cmb_d21_0.l_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13660\,
            in2 => \N__13843\,
            in3 => \N__12729\,
            lcout => \inst_midgetv_core.inst_shiftcounter.genblk1_d_0\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_shiftcounter.genblk1_reg_shcnt40_1_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__11998\,
            in1 => \N__11992\,
            in2 => \N__12539\,
            in3 => \N__11986\,
            lcout => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_1\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_0\,
            carryout => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_1\,
            clk => \N__13818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_shiftcounter.genblk1_reg_shcnt40_2_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__13636\,
            in1 => \N__12530\,
            in2 => \N__11983\,
            in3 => \N__11974\,
            lcout => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_2\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_1\,
            carryout => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_2\,
            clk => \N__13818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_shiftcounter.genblk1_reg_shcnt40_3_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__12757\,
            in1 => \N__13033\,
            in2 => \N__12540\,
            in3 => \N__13027\,
            lcout => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_3\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_2\,
            carryout => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_3\,
            clk => \N__13818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_shiftcounter.genblk1_reg_shcnt40_4_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__12664\,
            in1 => \N__12534\,
            in2 => \N__13024\,
            in3 => \N__13015\,
            lcout => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_4\,
            ltout => OPEN,
            carryin => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_3\,
            carryout => \inst_midgetv_core.inst_shiftcounter.genblk1_shcy_4\,
            clk => \N__13818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_shiftcounter.genblk1_cmb_lastshift.l_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__12535\,
            in1 => \N__12998\,
            in2 => \N__13010\,
            in3 => \N__12796\,
            lcout => \inst_midgetv_core.lastshift\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_shiftcounter.genblk1_cmb_d43_0.l_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__13668\,
            in1 => \N__14047\,
            in2 => \_gnd_net_\,
            in3 => \N__12477\,
            lcout => \inst_midgetv_core.inst_shiftcounter.genblk1_d_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_shiftcounter.genblk1_cmb_d43_1.l_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12728\,
            in1 => \N__13669\,
            in2 => \_gnd_net_\,
            in3 => \N__15127\,
            lcout => \inst_midgetv_core.inst_shiftcounter.genblk1_d_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.we_I_0_2_lut_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__12585\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12658\,
            lcout => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrb.we\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.we_I_0_2_lut_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__12586\,
            in1 => \_gnd_net_\,
            in2 => \N__12628\,
            in3 => \_gnd_net_\,
            lcout => \inst_midgetv_core.inst_ebr.ebrh.genblk1_ebrh.we\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.we_I_0_2_lut_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12595\,
            in2 => \_gnd_net_\,
            in3 => \N__12584\,
            lcout => \inst_midgetv_core.inst_ebr.ebrb.genblk1_ebrh.we\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_shiftcounter.genblk1_reg_shcnt40_0_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001001110010000"
        )
    port map (
            in0 => \N__13842\,
            in1 => \N__13667\,
            in2 => \N__12541\,
            in3 => \N__12499\,
            lcout => \inst_midgetv_core.inst_shiftcounter.dbg_rshcnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_shiftcounter.genblk1_cmb_d21_1.l_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__13666\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14194\,
            lcout => \inst_midgetv_core.inst_shiftcounter.genblk1_d_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_sel_3_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__13569\,
            in1 => \N__13585\,
            in2 => \N__13630\,
            in3 => \N__13536\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_sel_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_sel0hack_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__13583\,
            in1 => \N__13596\,
            in2 => \_gnd_net_\,
            in3 => \N__13608\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_sel0hack\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_sel0h_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011001"
        )
    port map (
            in0 => \N__13597\,
            in1 => \N__13584\,
            in2 => \N__13570\,
            in3 => \N__13535\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_sel0h\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_sel_0_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__13477\,
            in1 => \N__13462\,
            in2 => \_gnd_net_\,
            in3 => \N__13456\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_sel_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_wai.genblk1_L_2326_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__13450\,
            in1 => \_gnd_net_\,
            in2 => \N__13366\,
            in3 => \N__13273\,
            lcout => \inst_midgetv_core.Wai_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_b1a_LC_18_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__14569\,
            in1 => \N__14652\,
            in2 => \N__13180\,
            in3 => \N__13137\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_b1a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_b3a_LC_18_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__14570\,
            in1 => \N__14653\,
            in2 => \N__13105\,
            in3 => \N__13060\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_b3a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_ss1_LC_18_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15324\,
            in1 => \N__14007\,
            in2 => \_gnd_net_\,
            in3 => \N__15078\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_ss1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_b4a_LC_18_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__14654\,
            in1 => \N__14572\,
            in2 => \N__14472\,
            in3 => \N__14431\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_b4a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_ss0_LC_18_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15077\,
            in1 => \N__15323\,
            in2 => \_gnd_net_\,
            in3 => \N__14136\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_ss0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_b0a_LC_18_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__14651\,
            in1 => \N__14571\,
            in2 => \N__14395\,
            in3 => \N__14335\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_b0a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_Rai4_LC_18_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__14696\,
            in1 => \N__14302\,
            in2 => \_gnd_net_\,
            in3 => \N__14257\,
            lcout => \inst_midgetv_core.Rai_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_Rai0_LC_18_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001100"
        )
    port map (
            in0 => \N__14199\,
            in1 => \N__14137\,
            in2 => \N__14702\,
            in3 => \N__14119\,
            lcout => \inst_midgetv_core.Rai_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_Rai1_LC_18_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__14692\,
            in1 => \N__14062\,
            in2 => \N__14014\,
            in3 => \N__13984\,
            lcout => \inst_midgetv_core.Rai_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_Rai5_LC_18_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__14576\,
            in1 => \N__13926\,
            in2 => \_gnd_net_\,
            in3 => \N__14697\,
            lcout => \inst_midgetv_core.Rai_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_Rai3_LC_18_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001010"
        )
    port map (
            in0 => \N__15325\,
            in1 => \N__15307\,
            in2 => \N__14703\,
            in3 => \N__15262\,
            lcout => \inst_midgetv_core.Rai_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_b2a_LC_18_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__14682\,
            in1 => \N__14577\,
            in2 => \N__15205\,
            in3 => \N__15166\,
            lcout => \inst_midgetv_core.inst_rai.genblk1_b2a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_Rai2_LC_18_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__14683\,
            in1 => \N__15132\,
            in2 => \N__15082\,
            in3 => \N__15049\,
            lcout => \inst_midgetv_core.Rai_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_genblk1_L_Rai8_LC_18_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14684\,
            in1 => \N__14578\,
            in2 => \_gnd_net_\,
            in3 => \N__14992\,
            lcout => \inst_midgetv_core.Rai_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_genblk1_genblk1_L_Rai9_LC_18_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14685\,
            in1 => \N__14579\,
            in2 => \_gnd_net_\,
            in3 => \N__14892\,
            lcout => \inst_midgetv_core.Rai_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_Rai6_LC_20_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14704\,
            in1 => \N__14797\,
            in2 => \_gnd_net_\,
            in3 => \N__14587\,
            lcout => \inst_midgetv_core.Rai_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \inst_midgetv_core.inst_rai.genblk1_L_Rai7_LC_20_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14701\,
            in1 => \N__14619\,
            in2 => \_gnd_net_\,
            in3 => \N__14586\,
            lcout => \inst_midgetv_core.Rai_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
