/* -----------------------------------------------------------------------------
 * Part of midgetv
 * 2019. Copyright B. Nossum.
 * For licence, see LICENCE
 * -----------------------------------------------------------------------------
 * EBR holds constants, registers, and code. This is a wrapper,
 * EBRADRWIDTH  EBRs  Organization   Gives     Capacity  WRITE/READ mode
 *  8           2     16 x  8 *  2   32 x  8   1 kiB     0
 *  9           4      8 x  9 *  4   32 x  9   2 kiB     1
 * 10           8      4 x 10 *  8   32 x 10   4 kiB     2
 * 11           16     2 x 11 * 16   32 x 11   8 kiB     3
 * 
 * In this illustration, for brevity; m0 = bmask0 etc, w=iwe
 * EBRADRWIDTH
 *    EBR15 EBR14 EBR13 EBR12 EBR11 EBR10 EBR9  EBR8  EBR7  EBR6  EBR5  EBR4  EBR3  EBR2  EBR1  EBR0
 *  8                                                                                     w     w
 *  9                                                                         w&m3  w&m2  w&m1  w&m0
 * 10                                                 w&m3  w&m3  w&m2  w&m2  w&m1  w&m1  w&m0  w&m0
 * 11 w&m3  w&m3  w&m3  w&m3  ie&m2 ie&m2 ie&m2 ie&m2 w&m1  w&m1  w&m1  w&m1  w&m0  w&m0  w&m0  w&m0
 * 
 */
module m_ebr
  # ( parameter EBRADRWIDTH = 8,
      parameter [4095:0] prg00 = 4096'h0,
      parameter [4095:0] prg01 = 4096'h0,
      parameter [4095:0] prg02 = 4096'h0,
      parameter [4095:0] prg03 = 4096'h0,
      parameter [4095:0] prg04 = 4096'h0,
      parameter [4095:0] prg05 = 4096'h0,
      parameter [4095:0] prg06 = 4096'h0,
      parameter [4095:0] prg07 = 4096'h0,
      parameter [4095:0] prg08 = 4096'h0,
      parameter [4095:0] prg09 = 4096'h0,
      parameter [4095:0] prg0A = 4096'h0,
      parameter [4095:0] prg0B = 4096'h0,
      parameter [4095:0] prg0C = 4096'h0,
      parameter [4095:0] prg0D = 4096'h0,
      parameter [4095:0] prg0E = 4096'h0,
      parameter [4095:0] prg0F = 4096'h0
      )
   (
    input [31:0]            B, //     Output from ALU
    input [EBRADRWIDTH-1:0] Rai, //   Read address
    input [EBRADRWIDTH-1:0] Wai, //   Write address    
    input                   clk, //   System clock
    input [3:0]             bmask, // Byte masks for write, active LOW
    input                   iwe, //   Write enable
    output [31:0]           DAT_O, //  Register used in many places, also I/O output
    output                  next_readvalue_unknown // For debugging only
    );
   wire [31:0]              eDAT_O;
`ifdef verilator 
   reg                      readvalue_unknown;
   assign next_readvalue_unknown =  ( Rai == Wai && iwe );
   always @(posedge clk)
     readvalue_unknown <= next_readvalue_unknown;
   assign DAT_O = readvalue_unknown ? 32'hdeaddead : eDAT_O;
`else
   assign next_readvalue_unknown = 1'b0;
   assign DAT_O = eDAT_O;
`endif

   /* Split the up to 8 KiB program into low and high halfword
    */
   localparam [4095:0]
     pb7 = {prg0F[4079:4064],prg0F[4047:4032],prg0F[4015:4000],prg0F[3983:3968],prg0F[3951:3936],prg0F[3919:3904],prg0F[3887:3872],prg0F[3855:3840],
            prg0F[3823:3808],prg0F[3791:3776],prg0F[3759:3744],prg0F[3727:3712],prg0F[3695:3680],prg0F[3663:3648],prg0F[3631:3616],prg0F[3599:3584],
            prg0F[3567:3552],prg0F[3535:3520],prg0F[3503:3488],prg0F[3471:3456],prg0F[3439:3424],prg0F[3407:3392],prg0F[3375:3360],prg0F[3343:3328],
            prg0F[3311:3296],prg0F[3279:3264],prg0F[3247:3232],prg0F[3215:3200],prg0F[3183:3168],prg0F[3151:3136],prg0F[3119:3104],prg0F[3087:3072],
            prg0F[3055:3040],prg0F[3023:3008],prg0F[2991:2976],prg0F[2959:2944],prg0F[2927:2912],prg0F[2895:2880],prg0F[2863:2848],prg0F[2831:2816],
            prg0F[2799:2784],prg0F[2767:2752],prg0F[2735:2720],prg0F[2703:2688],prg0F[2671:2656],prg0F[2639:2624],prg0F[2607:2592],prg0F[2575:2560],
            prg0F[2543:2528],prg0F[2511:2496],prg0F[2479:2464],prg0F[2447:2432],prg0F[2415:2400],prg0F[2383:2368],prg0F[2351:2336],prg0F[2319:2304],
            prg0F[2287:2272],prg0F[2255:2240],prg0F[2223:2208],prg0F[2191:2176],prg0F[2159:2144],prg0F[2127:2112],prg0F[2095:2080],prg0F[2063:2048],
            prg0F[2031:2016],prg0F[1999:1984],prg0F[1967:1952],prg0F[1935:1920],prg0F[1903:1888],prg0F[1871:1856],prg0F[1839:1824],prg0F[1807:1792],
            prg0F[1775:1760],prg0F[1743:1728],prg0F[1711:1696],prg0F[1679:1664],prg0F[1647:1632],prg0F[1615:1600],prg0F[1583:1568],prg0F[1551:1536],
            prg0F[1519:1504],prg0F[1487:1472],prg0F[1455:1440],prg0F[1423:1408],prg0F[1391:1376],prg0F[1359:1344],prg0F[1327:1312],prg0F[1295:1280],
            prg0F[1263:1248],prg0F[1231:1216],prg0F[1199:1184],prg0F[1167:1152],prg0F[1135:1120],prg0F[1103:1088],prg0F[1071:1056],prg0F[1039:1024],
            prg0F[1007: 992],prg0F[ 975: 960],prg0F[ 943: 928],prg0F[ 911: 896],prg0F[ 879: 864],prg0F[ 847: 832],prg0F[ 815: 800],prg0F[ 783: 768],
            prg0F[ 751: 736],prg0F[ 719: 704],prg0F[ 687: 672],prg0F[ 655: 640],prg0F[ 623: 608],prg0F[ 591: 576],prg0F[ 559: 544],prg0F[ 527: 512],
            prg0F[ 495: 480],prg0F[ 463: 448],prg0F[ 431: 416],prg0F[ 399: 384],prg0F[ 367: 352],prg0F[ 335: 320],prg0F[ 303: 288],prg0F[ 271: 256],
            prg0F[ 239: 224],prg0F[ 207: 192],prg0F[ 175: 160],prg0F[ 143: 128],prg0F[ 111:  96],prg0F[  79:  64],prg0F[  47:  32],prg0F[  15:   0],
            prg0E[4079:4064],prg0E[4047:4032],prg0E[4015:4000],prg0E[3983:3968],prg0E[3951:3936],prg0E[3919:3904],prg0E[3887:3872],prg0E[3855:3840],
            prg0E[3823:3808],prg0E[3791:3776],prg0E[3759:3744],prg0E[3727:3712],prg0E[3695:3680],prg0E[3663:3648],prg0E[3631:3616],prg0E[3599:3584],
            prg0E[3567:3552],prg0E[3535:3520],prg0E[3503:3488],prg0E[3471:3456],prg0E[3439:3424],prg0E[3407:3392],prg0E[3375:3360],prg0E[3343:3328],
            prg0E[3311:3296],prg0E[3279:3264],prg0E[3247:3232],prg0E[3215:3200],prg0E[3183:3168],prg0E[3151:3136],prg0E[3119:3104],prg0E[3087:3072],
            prg0E[3055:3040],prg0E[3023:3008],prg0E[2991:2976],prg0E[2959:2944],prg0E[2927:2912],prg0E[2895:2880],prg0E[2863:2848],prg0E[2831:2816],
            prg0E[2799:2784],prg0E[2767:2752],prg0E[2735:2720],prg0E[2703:2688],prg0E[2671:2656],prg0E[2639:2624],prg0E[2607:2592],prg0E[2575:2560],
            prg0E[2543:2528],prg0E[2511:2496],prg0E[2479:2464],prg0E[2447:2432],prg0E[2415:2400],prg0E[2383:2368],prg0E[2351:2336],prg0E[2319:2304],
            prg0E[2287:2272],prg0E[2255:2240],prg0E[2223:2208],prg0E[2191:2176],prg0E[2159:2144],prg0E[2127:2112],prg0E[2095:2080],prg0E[2063:2048],
            prg0E[2031:2016],prg0E[1999:1984],prg0E[1967:1952],prg0E[1935:1920],prg0E[1903:1888],prg0E[1871:1856],prg0E[1839:1824],prg0E[1807:1792],
            prg0E[1775:1760],prg0E[1743:1728],prg0E[1711:1696],prg0E[1679:1664],prg0E[1647:1632],prg0E[1615:1600],prg0E[1583:1568],prg0E[1551:1536],
            prg0E[1519:1504],prg0E[1487:1472],prg0E[1455:1440],prg0E[1423:1408],prg0E[1391:1376],prg0E[1359:1344],prg0E[1327:1312],prg0E[1295:1280],
            prg0E[1263:1248],prg0E[1231:1216],prg0E[1199:1184],prg0E[1167:1152],prg0E[1135:1120],prg0E[1103:1088],prg0E[1071:1056],prg0E[1039:1024],
            prg0E[1007: 992],prg0E[ 975: 960],prg0E[ 943: 928],prg0E[ 911: 896],prg0E[ 879: 864],prg0E[ 847: 832],prg0E[ 815: 800],prg0E[ 783: 768],
            prg0E[ 751: 736],prg0E[ 719: 704],prg0E[ 687: 672],prg0E[ 655: 640],prg0E[ 623: 608],prg0E[ 591: 576],prg0E[ 559: 544],prg0E[ 527: 512],
            prg0E[ 495: 480],prg0E[ 463: 448],prg0E[ 431: 416],prg0E[ 399: 384],prg0E[ 367: 352],prg0E[ 335: 320],prg0E[ 303: 288],prg0E[ 271: 256],
            prg0E[ 239: 224],prg0E[ 207: 192],prg0E[ 175: 160],prg0E[ 143: 128],prg0E[ 111:  96],prg0E[  79:  64],prg0E[  47:  32],prg0E[  15:   0]};
   localparam [4095:0]
     pb6 = {prg0D[4079:4064],prg0D[4047:4032],prg0D[4015:4000],prg0D[3983:3968],prg0D[3951:3936],prg0D[3919:3904],prg0D[3887:3872],prg0D[3855:3840],
            prg0D[3823:3808],prg0D[3791:3776],prg0D[3759:3744],prg0D[3727:3712],prg0D[3695:3680],prg0D[3663:3648],prg0D[3631:3616],prg0D[3599:3584],
            prg0D[3567:3552],prg0D[3535:3520],prg0D[3503:3488],prg0D[3471:3456],prg0D[3439:3424],prg0D[3407:3392],prg0D[3375:3360],prg0D[3343:3328],
            prg0D[3311:3296],prg0D[3279:3264],prg0D[3247:3232],prg0D[3215:3200],prg0D[3183:3168],prg0D[3151:3136],prg0D[3119:3104],prg0D[3087:3072],
            prg0D[3055:3040],prg0D[3023:3008],prg0D[2991:2976],prg0D[2959:2944],prg0D[2927:2912],prg0D[2895:2880],prg0D[2863:2848],prg0D[2831:2816],
            prg0D[2799:2784],prg0D[2767:2752],prg0D[2735:2720],prg0D[2703:2688],prg0D[2671:2656],prg0D[2639:2624],prg0D[2607:2592],prg0D[2575:2560],
            prg0D[2543:2528],prg0D[2511:2496],prg0D[2479:2464],prg0D[2447:2432],prg0D[2415:2400],prg0D[2383:2368],prg0D[2351:2336],prg0D[2319:2304],
            prg0D[2287:2272],prg0D[2255:2240],prg0D[2223:2208],prg0D[2191:2176],prg0D[2159:2144],prg0D[2127:2112],prg0D[2095:2080],prg0D[2063:2048],
            prg0D[2031:2016],prg0D[1999:1984],prg0D[1967:1952],prg0D[1935:1920],prg0D[1903:1888],prg0D[1871:1856],prg0D[1839:1824],prg0D[1807:1792],
            prg0D[1775:1760],prg0D[1743:1728],prg0D[1711:1696],prg0D[1679:1664],prg0D[1647:1632],prg0D[1615:1600],prg0D[1583:1568],prg0D[1551:1536],
            prg0D[1519:1504],prg0D[1487:1472],prg0D[1455:1440],prg0D[1423:1408],prg0D[1391:1376],prg0D[1359:1344],prg0D[1327:1312],prg0D[1295:1280],
            prg0D[1263:1248],prg0D[1231:1216],prg0D[1199:1184],prg0D[1167:1152],prg0D[1135:1120],prg0D[1103:1088],prg0D[1071:1056],prg0D[1039:1024],
            prg0D[1007: 992],prg0D[ 975: 960],prg0D[ 943: 928],prg0D[ 911: 896],prg0D[ 879: 864],prg0D[ 847: 832],prg0D[ 815: 800],prg0D[ 783: 768],
            prg0D[ 751: 736],prg0D[ 719: 704],prg0D[ 687: 672],prg0D[ 655: 640],prg0D[ 623: 608],prg0D[ 591: 576],prg0D[ 559: 544],prg0D[ 527: 512],
            prg0D[ 495: 480],prg0D[ 463: 448],prg0D[ 431: 416],prg0D[ 399: 384],prg0D[ 367: 352],prg0D[ 335: 320],prg0D[ 303: 288],prg0D[ 271: 256],
            prg0D[ 239: 224],prg0D[ 207: 192],prg0D[ 175: 160],prg0D[ 143: 128],prg0D[ 111:  96],prg0D[  79:  64],prg0D[  47:  32],prg0D[  15:   0],
            prg0C[4079:4064],prg0C[4047:4032],prg0C[4015:4000],prg0C[3983:3968],prg0C[3951:3936],prg0C[3919:3904],prg0C[3887:3872],prg0C[3855:3840],
            prg0C[3823:3808],prg0C[3791:3776],prg0C[3759:3744],prg0C[3727:3712],prg0C[3695:3680],prg0C[3663:3648],prg0C[3631:3616],prg0C[3599:3584],
            prg0C[3567:3552],prg0C[3535:3520],prg0C[3503:3488],prg0C[3471:3456],prg0C[3439:3424],prg0C[3407:3392],prg0C[3375:3360],prg0C[3343:3328],
            prg0C[3311:3296],prg0C[3279:3264],prg0C[3247:3232],prg0C[3215:3200],prg0C[3183:3168],prg0C[3151:3136],prg0C[3119:3104],prg0C[3087:3072],
            prg0C[3055:3040],prg0C[3023:3008],prg0C[2991:2976],prg0C[2959:2944],prg0C[2927:2912],prg0C[2895:2880],prg0C[2863:2848],prg0C[2831:2816],
            prg0C[2799:2784],prg0C[2767:2752],prg0C[2735:2720],prg0C[2703:2688],prg0C[2671:2656],prg0C[2639:2624],prg0C[2607:2592],prg0C[2575:2560],
            prg0C[2543:2528],prg0C[2511:2496],prg0C[2479:2464],prg0C[2447:2432],prg0C[2415:2400],prg0C[2383:2368],prg0C[2351:2336],prg0C[2319:2304],
            prg0C[2287:2272],prg0C[2255:2240],prg0C[2223:2208],prg0C[2191:2176],prg0C[2159:2144],prg0C[2127:2112],prg0C[2095:2080],prg0C[2063:2048],
            prg0C[2031:2016],prg0C[1999:1984],prg0C[1967:1952],prg0C[1935:1920],prg0C[1903:1888],prg0C[1871:1856],prg0C[1839:1824],prg0C[1807:1792],
            prg0C[1775:1760],prg0C[1743:1728],prg0C[1711:1696],prg0C[1679:1664],prg0C[1647:1632],prg0C[1615:1600],prg0C[1583:1568],prg0C[1551:1536],
            prg0C[1519:1504],prg0C[1487:1472],prg0C[1455:1440],prg0C[1423:1408],prg0C[1391:1376],prg0C[1359:1344],prg0C[1327:1312],prg0C[1295:1280],
            prg0C[1263:1248],prg0C[1231:1216],prg0C[1199:1184],prg0C[1167:1152],prg0C[1135:1120],prg0C[1103:1088],prg0C[1071:1056],prg0C[1039:1024],
            prg0C[1007: 992],prg0C[ 975: 960],prg0C[ 943: 928],prg0C[ 911: 896],prg0C[ 879: 864],prg0C[ 847: 832],prg0C[ 815: 800],prg0C[ 783: 768],
            prg0C[ 751: 736],prg0C[ 719: 704],prg0C[ 687: 672],prg0C[ 655: 640],prg0C[ 623: 608],prg0C[ 591: 576],prg0C[ 559: 544],prg0C[ 527: 512],
            prg0C[ 495: 480],prg0C[ 463: 448],prg0C[ 431: 416],prg0C[ 399: 384],prg0C[ 367: 352],prg0C[ 335: 320],prg0C[ 303: 288],prg0C[ 271: 256],
            prg0C[ 239: 224],prg0C[ 207: 192],prg0C[ 175: 160],prg0C[ 143: 128],prg0C[ 111:  96],prg0C[  79:  64],prg0C[  47:  32],prg0C[  15:   0]};
   localparam [4095:0]
     pb5 = {prg0B[4079:4064],prg0B[4047:4032],prg0B[4015:4000],prg0B[3983:3968],prg0B[3951:3936],prg0B[3919:3904],prg0B[3887:3872],prg0B[3855:3840],
            prg0B[3823:3808],prg0B[3791:3776],prg0B[3759:3744],prg0B[3727:3712],prg0B[3695:3680],prg0B[3663:3648],prg0B[3631:3616],prg0B[3599:3584],
            prg0B[3567:3552],prg0B[3535:3520],prg0B[3503:3488],prg0B[3471:3456],prg0B[3439:3424],prg0B[3407:3392],prg0B[3375:3360],prg0B[3343:3328],
            prg0B[3311:3296],prg0B[3279:3264],prg0B[3247:3232],prg0B[3215:3200],prg0B[3183:3168],prg0B[3151:3136],prg0B[3119:3104],prg0B[3087:3072],
            prg0B[3055:3040],prg0B[3023:3008],prg0B[2991:2976],prg0B[2959:2944],prg0B[2927:2912],prg0B[2895:2880],prg0B[2863:2848],prg0B[2831:2816],
            prg0B[2799:2784],prg0B[2767:2752],prg0B[2735:2720],prg0B[2703:2688],prg0B[2671:2656],prg0B[2639:2624],prg0B[2607:2592],prg0B[2575:2560],
            prg0B[2543:2528],prg0B[2511:2496],prg0B[2479:2464],prg0B[2447:2432],prg0B[2415:2400],prg0B[2383:2368],prg0B[2351:2336],prg0B[2319:2304],
            prg0B[2287:2272],prg0B[2255:2240],prg0B[2223:2208],prg0B[2191:2176],prg0B[2159:2144],prg0B[2127:2112],prg0B[2095:2080],prg0B[2063:2048],
            prg0B[2031:2016],prg0B[1999:1984],prg0B[1967:1952],prg0B[1935:1920],prg0B[1903:1888],prg0B[1871:1856],prg0B[1839:1824],prg0B[1807:1792],
            prg0B[1775:1760],prg0B[1743:1728],prg0B[1711:1696],prg0B[1679:1664],prg0B[1647:1632],prg0B[1615:1600],prg0B[1583:1568],prg0B[1551:1536],
            prg0B[1519:1504],prg0B[1487:1472],prg0B[1455:1440],prg0B[1423:1408],prg0B[1391:1376],prg0B[1359:1344],prg0B[1327:1312],prg0B[1295:1280],
            prg0B[1263:1248],prg0B[1231:1216],prg0B[1199:1184],prg0B[1167:1152],prg0B[1135:1120],prg0B[1103:1088],prg0B[1071:1056],prg0B[1039:1024],
            prg0B[1007: 992],prg0B[ 975: 960],prg0B[ 943: 928],prg0B[ 911: 896],prg0B[ 879: 864],prg0B[ 847: 832],prg0B[ 815: 800],prg0B[ 783: 768],
            prg0B[ 751: 736],prg0B[ 719: 704],prg0B[ 687: 672],prg0B[ 655: 640],prg0B[ 623: 608],prg0B[ 591: 576],prg0B[ 559: 544],prg0B[ 527: 512],
            prg0B[ 495: 480],prg0B[ 463: 448],prg0B[ 431: 416],prg0B[ 399: 384],prg0B[ 367: 352],prg0B[ 335: 320],prg0B[ 303: 288],prg0B[ 271: 256],
            prg0B[ 239: 224],prg0B[ 207: 192],prg0B[ 175: 160],prg0B[ 143: 128],prg0B[ 111:  96],prg0B[  79:  64],prg0B[  47:  32],prg0B[  15:   0],
            prg0A[4079:4064],prg0A[4047:4032],prg0A[4015:4000],prg0A[3983:3968],prg0A[3951:3936],prg0A[3919:3904],prg0A[3887:3872],prg0A[3855:3840],
            prg0A[3823:3808],prg0A[3791:3776],prg0A[3759:3744],prg0A[3727:3712],prg0A[3695:3680],prg0A[3663:3648],prg0A[3631:3616],prg0A[3599:3584],
            prg0A[3567:3552],prg0A[3535:3520],prg0A[3503:3488],prg0A[3471:3456],prg0A[3439:3424],prg0A[3407:3392],prg0A[3375:3360],prg0A[3343:3328],
            prg0A[3311:3296],prg0A[3279:3264],prg0A[3247:3232],prg0A[3215:3200],prg0A[3183:3168],prg0A[3151:3136],prg0A[3119:3104],prg0A[3087:3072],
            prg0A[3055:3040],prg0A[3023:3008],prg0A[2991:2976],prg0A[2959:2944],prg0A[2927:2912],prg0A[2895:2880],prg0A[2863:2848],prg0A[2831:2816],
            prg0A[2799:2784],prg0A[2767:2752],prg0A[2735:2720],prg0A[2703:2688],prg0A[2671:2656],prg0A[2639:2624],prg0A[2607:2592],prg0A[2575:2560],
            prg0A[2543:2528],prg0A[2511:2496],prg0A[2479:2464],prg0A[2447:2432],prg0A[2415:2400],prg0A[2383:2368],prg0A[2351:2336],prg0A[2319:2304],
            prg0A[2287:2272],prg0A[2255:2240],prg0A[2223:2208],prg0A[2191:2176],prg0A[2159:2144],prg0A[2127:2112],prg0A[2095:2080],prg0A[2063:2048],
            prg0A[2031:2016],prg0A[1999:1984],prg0A[1967:1952],prg0A[1935:1920],prg0A[1903:1888],prg0A[1871:1856],prg0A[1839:1824],prg0A[1807:1792],
            prg0A[1775:1760],prg0A[1743:1728],prg0A[1711:1696],prg0A[1679:1664],prg0A[1647:1632],prg0A[1615:1600],prg0A[1583:1568],prg0A[1551:1536],
            prg0A[1519:1504],prg0A[1487:1472],prg0A[1455:1440],prg0A[1423:1408],prg0A[1391:1376],prg0A[1359:1344],prg0A[1327:1312],prg0A[1295:1280],
            prg0A[1263:1248],prg0A[1231:1216],prg0A[1199:1184],prg0A[1167:1152],prg0A[1135:1120],prg0A[1103:1088],prg0A[1071:1056],prg0A[1039:1024],
            prg0A[1007: 992],prg0A[ 975: 960],prg0A[ 943: 928],prg0A[ 911: 896],prg0A[ 879: 864],prg0A[ 847: 832],prg0A[ 815: 800],prg0A[ 783: 768],
            prg0A[ 751: 736],prg0A[ 719: 704],prg0A[ 687: 672],prg0A[ 655: 640],prg0A[ 623: 608],prg0A[ 591: 576],prg0A[ 559: 544],prg0A[ 527: 512],
            prg0A[ 495: 480],prg0A[ 463: 448],prg0A[ 431: 416],prg0A[ 399: 384],prg0A[ 367: 352],prg0A[ 335: 320],prg0A[ 303: 288],prg0A[ 271: 256],
            prg0A[ 239: 224],prg0A[ 207: 192],prg0A[ 175: 160],prg0A[ 143: 128],prg0A[ 111:  96],prg0A[  79:  64],prg0A[  47:  32],prg0A[  15:   0]};
   localparam [4095:0]
     pb4 = {prg09[4079:4064],prg09[4047:4032],prg09[4015:4000],prg09[3983:3968],prg09[3951:3936],prg09[3919:3904],prg09[3887:3872],prg09[3855:3840],
            prg09[3823:3808],prg09[3791:3776],prg09[3759:3744],prg09[3727:3712],prg09[3695:3680],prg09[3663:3648],prg09[3631:3616],prg09[3599:3584],
            prg09[3567:3552],prg09[3535:3520],prg09[3503:3488],prg09[3471:3456],prg09[3439:3424],prg09[3407:3392],prg09[3375:3360],prg09[3343:3328],
            prg09[3311:3296],prg09[3279:3264],prg09[3247:3232],prg09[3215:3200],prg09[3183:3168],prg09[3151:3136],prg09[3119:3104],prg09[3087:3072],
            prg09[3055:3040],prg09[3023:3008],prg09[2991:2976],prg09[2959:2944],prg09[2927:2912],prg09[2895:2880],prg09[2863:2848],prg09[2831:2816],
            prg09[2799:2784],prg09[2767:2752],prg09[2735:2720],prg09[2703:2688],prg09[2671:2656],prg09[2639:2624],prg09[2607:2592],prg09[2575:2560],
            prg09[2543:2528],prg09[2511:2496],prg09[2479:2464],prg09[2447:2432],prg09[2415:2400],prg09[2383:2368],prg09[2351:2336],prg09[2319:2304],
            prg09[2287:2272],prg09[2255:2240],prg09[2223:2208],prg09[2191:2176],prg09[2159:2144],prg09[2127:2112],prg09[2095:2080],prg09[2063:2048],
            prg09[2031:2016],prg09[1999:1984],prg09[1967:1952],prg09[1935:1920],prg09[1903:1888],prg09[1871:1856],prg09[1839:1824],prg09[1807:1792],
            prg09[1775:1760],prg09[1743:1728],prg09[1711:1696],prg09[1679:1664],prg09[1647:1632],prg09[1615:1600],prg09[1583:1568],prg09[1551:1536],
            prg09[1519:1504],prg09[1487:1472],prg09[1455:1440],prg09[1423:1408],prg09[1391:1376],prg09[1359:1344],prg09[1327:1312],prg09[1295:1280],
            prg09[1263:1248],prg09[1231:1216],prg09[1199:1184],prg09[1167:1152],prg09[1135:1120],prg09[1103:1088],prg09[1071:1056],prg09[1039:1024],
            prg09[1007: 992],prg09[ 975: 960],prg09[ 943: 928],prg09[ 911: 896],prg09[ 879: 864],prg09[ 847: 832],prg09[ 815: 800],prg09[ 783: 768],
            prg09[ 751: 736],prg09[ 719: 704],prg09[ 687: 672],prg09[ 655: 640],prg09[ 623: 608],prg09[ 591: 576],prg09[ 559: 544],prg09[ 527: 512],
            prg09[ 495: 480],prg09[ 463: 448],prg09[ 431: 416],prg09[ 399: 384],prg09[ 367: 352],prg09[ 335: 320],prg09[ 303: 288],prg09[ 271: 256],
            prg09[ 239: 224],prg09[ 207: 192],prg09[ 175: 160],prg09[ 143: 128],prg09[ 111:  96],prg09[  79:  64],prg09[  47:  32],prg09[  15:   0],
            prg08[4079:4064],prg08[4047:4032],prg08[4015:4000],prg08[3983:3968],prg08[3951:3936],prg08[3919:3904],prg08[3887:3872],prg08[3855:3840],
            prg08[3823:3808],prg08[3791:3776],prg08[3759:3744],prg08[3727:3712],prg08[3695:3680],prg08[3663:3648],prg08[3631:3616],prg08[3599:3584],
            prg08[3567:3552],prg08[3535:3520],prg08[3503:3488],prg08[3471:3456],prg08[3439:3424],prg08[3407:3392],prg08[3375:3360],prg08[3343:3328],
            prg08[3311:3296],prg08[3279:3264],prg08[3247:3232],prg08[3215:3200],prg08[3183:3168],prg08[3151:3136],prg08[3119:3104],prg08[3087:3072],
            prg08[3055:3040],prg08[3023:3008],prg08[2991:2976],prg08[2959:2944],prg08[2927:2912],prg08[2895:2880],prg08[2863:2848],prg08[2831:2816],
            prg08[2799:2784],prg08[2767:2752],prg08[2735:2720],prg08[2703:2688],prg08[2671:2656],prg08[2639:2624],prg08[2607:2592],prg08[2575:2560],
            prg08[2543:2528],prg08[2511:2496],prg08[2479:2464],prg08[2447:2432],prg08[2415:2400],prg08[2383:2368],prg08[2351:2336],prg08[2319:2304],
            prg08[2287:2272],prg08[2255:2240],prg08[2223:2208],prg08[2191:2176],prg08[2159:2144],prg08[2127:2112],prg08[2095:2080],prg08[2063:2048],
            prg08[2031:2016],prg08[1999:1984],prg08[1967:1952],prg08[1935:1920],prg08[1903:1888],prg08[1871:1856],prg08[1839:1824],prg08[1807:1792],
            prg08[1775:1760],prg08[1743:1728],prg08[1711:1696],prg08[1679:1664],prg08[1647:1632],prg08[1615:1600],prg08[1583:1568],prg08[1551:1536],
            prg08[1519:1504],prg08[1487:1472],prg08[1455:1440],prg08[1423:1408],prg08[1391:1376],prg08[1359:1344],prg08[1327:1312],prg08[1295:1280],
            prg08[1263:1248],prg08[1231:1216],prg08[1199:1184],prg08[1167:1152],prg08[1135:1120],prg08[1103:1088],prg08[1071:1056],prg08[1039:1024],
            prg08[1007: 992],prg08[ 975: 960],prg08[ 943: 928],prg08[ 911: 896],prg08[ 879: 864],prg08[ 847: 832],prg08[ 815: 800],prg08[ 783: 768],
            prg08[ 751: 736],prg08[ 719: 704],prg08[ 687: 672],prg08[ 655: 640],prg08[ 623: 608],prg08[ 591: 576],prg08[ 559: 544],prg08[ 527: 512],
            prg08[ 495: 480],prg08[ 463: 448],prg08[ 431: 416],prg08[ 399: 384],prg08[ 367: 352],prg08[ 335: 320],prg08[ 303: 288],prg08[ 271: 256],
            prg08[ 239: 224],prg08[ 207: 192],prg08[ 175: 160],prg08[ 143: 128],prg08[ 111:  96],prg08[  79:  64],prg08[  47:  32],prg08[  15:   0]};
   localparam [4095:0]
     pb3 = {prg07[4079:4064],prg07[4047:4032],prg07[4015:4000],prg07[3983:3968],prg07[3951:3936],prg07[3919:3904],prg07[3887:3872],prg07[3855:3840],
            prg07[3823:3808],prg07[3791:3776],prg07[3759:3744],prg07[3727:3712],prg07[3695:3680],prg07[3663:3648],prg07[3631:3616],prg07[3599:3584],
            prg07[3567:3552],prg07[3535:3520],prg07[3503:3488],prg07[3471:3456],prg07[3439:3424],prg07[3407:3392],prg07[3375:3360],prg07[3343:3328],
            prg07[3311:3296],prg07[3279:3264],prg07[3247:3232],prg07[3215:3200],prg07[3183:3168],prg07[3151:3136],prg07[3119:3104],prg07[3087:3072],
            prg07[3055:3040],prg07[3023:3008],prg07[2991:2976],prg07[2959:2944],prg07[2927:2912],prg07[2895:2880],prg07[2863:2848],prg07[2831:2816],
            prg07[2799:2784],prg07[2767:2752],prg07[2735:2720],prg07[2703:2688],prg07[2671:2656],prg07[2639:2624],prg07[2607:2592],prg07[2575:2560],
            prg07[2543:2528],prg07[2511:2496],prg07[2479:2464],prg07[2447:2432],prg07[2415:2400],prg07[2383:2368],prg07[2351:2336],prg07[2319:2304],
            prg07[2287:2272],prg07[2255:2240],prg07[2223:2208],prg07[2191:2176],prg07[2159:2144],prg07[2127:2112],prg07[2095:2080],prg07[2063:2048],
            prg07[2031:2016],prg07[1999:1984],prg07[1967:1952],prg07[1935:1920],prg07[1903:1888],prg07[1871:1856],prg07[1839:1824],prg07[1807:1792],
            prg07[1775:1760],prg07[1743:1728],prg07[1711:1696],prg07[1679:1664],prg07[1647:1632],prg07[1615:1600],prg07[1583:1568],prg07[1551:1536],
            prg07[1519:1504],prg07[1487:1472],prg07[1455:1440],prg07[1423:1408],prg07[1391:1376],prg07[1359:1344],prg07[1327:1312],prg07[1295:1280],
            prg07[1263:1248],prg07[1231:1216],prg07[1199:1184],prg07[1167:1152],prg07[1135:1120],prg07[1103:1088],prg07[1071:1056],prg07[1039:1024],
            prg07[1007: 992],prg07[ 975: 960],prg07[ 943: 928],prg07[ 911: 896],prg07[ 879: 864],prg07[ 847: 832],prg07[ 815: 800],prg07[ 783: 768],
            prg07[ 751: 736],prg07[ 719: 704],prg07[ 687: 672],prg07[ 655: 640],prg07[ 623: 608],prg07[ 591: 576],prg07[ 559: 544],prg07[ 527: 512],
            prg07[ 495: 480],prg07[ 463: 448],prg07[ 431: 416],prg07[ 399: 384],prg07[ 367: 352],prg07[ 335: 320],prg07[ 303: 288],prg07[ 271: 256],
            prg07[ 239: 224],prg07[ 207: 192],prg07[ 175: 160],prg07[ 143: 128],prg07[ 111:  96],prg07[  79:  64],prg07[  47:  32],prg07[  15:   0],
            prg06[4079:4064],prg06[4047:4032],prg06[4015:4000],prg06[3983:3968],prg06[3951:3936],prg06[3919:3904],prg06[3887:3872],prg06[3855:3840],
            prg06[3823:3808],prg06[3791:3776],prg06[3759:3744],prg06[3727:3712],prg06[3695:3680],prg06[3663:3648],prg06[3631:3616],prg06[3599:3584],
            prg06[3567:3552],prg06[3535:3520],prg06[3503:3488],prg06[3471:3456],prg06[3439:3424],prg06[3407:3392],prg06[3375:3360],prg06[3343:3328],
            prg06[3311:3296],prg06[3279:3264],prg06[3247:3232],prg06[3215:3200],prg06[3183:3168],prg06[3151:3136],prg06[3119:3104],prg06[3087:3072],
            prg06[3055:3040],prg06[3023:3008],prg06[2991:2976],prg06[2959:2944],prg06[2927:2912],prg06[2895:2880],prg06[2863:2848],prg06[2831:2816],
            prg06[2799:2784],prg06[2767:2752],prg06[2735:2720],prg06[2703:2688],prg06[2671:2656],prg06[2639:2624],prg06[2607:2592],prg06[2575:2560],
            prg06[2543:2528],prg06[2511:2496],prg06[2479:2464],prg06[2447:2432],prg06[2415:2400],prg06[2383:2368],prg06[2351:2336],prg06[2319:2304],
            prg06[2287:2272],prg06[2255:2240],prg06[2223:2208],prg06[2191:2176],prg06[2159:2144],prg06[2127:2112],prg06[2095:2080],prg06[2063:2048],
            prg06[2031:2016],prg06[1999:1984],prg06[1967:1952],prg06[1935:1920],prg06[1903:1888],prg06[1871:1856],prg06[1839:1824],prg06[1807:1792],
            prg06[1775:1760],prg06[1743:1728],prg06[1711:1696],prg06[1679:1664],prg06[1647:1632],prg06[1615:1600],prg06[1583:1568],prg06[1551:1536],
            prg06[1519:1504],prg06[1487:1472],prg06[1455:1440],prg06[1423:1408],prg06[1391:1376],prg06[1359:1344],prg06[1327:1312],prg06[1295:1280],
            prg06[1263:1248],prg06[1231:1216],prg06[1199:1184],prg06[1167:1152],prg06[1135:1120],prg06[1103:1088],prg06[1071:1056],prg06[1039:1024],
            prg06[1007: 992],prg06[ 975: 960],prg06[ 943: 928],prg06[ 911: 896],prg06[ 879: 864],prg06[ 847: 832],prg06[ 815: 800],prg06[ 783: 768],
            prg06[ 751: 736],prg06[ 719: 704],prg06[ 687: 672],prg06[ 655: 640],prg06[ 623: 608],prg06[ 591: 576],prg06[ 559: 544],prg06[ 527: 512],
            prg06[ 495: 480],prg06[ 463: 448],prg06[ 431: 416],prg06[ 399: 384],prg06[ 367: 352],prg06[ 335: 320],prg06[ 303: 288],prg06[ 271: 256],
            prg06[ 239: 224],prg06[ 207: 192],prg06[ 175: 160],prg06[ 143: 128],prg06[ 111:  96],prg06[  79:  64],prg06[  47:  32],prg06[  15:   0]};
   localparam [4095:0]
     pb2 = {prg05[4079:4064],prg05[4047:4032],prg05[4015:4000],prg05[3983:3968],prg05[3951:3936],prg05[3919:3904],prg05[3887:3872],prg05[3855:3840],
            prg05[3823:3808],prg05[3791:3776],prg05[3759:3744],prg05[3727:3712],prg05[3695:3680],prg05[3663:3648],prg05[3631:3616],prg05[3599:3584],
            prg05[3567:3552],prg05[3535:3520],prg05[3503:3488],prg05[3471:3456],prg05[3439:3424],prg05[3407:3392],prg05[3375:3360],prg05[3343:3328],
            prg05[3311:3296],prg05[3279:3264],prg05[3247:3232],prg05[3215:3200],prg05[3183:3168],prg05[3151:3136],prg05[3119:3104],prg05[3087:3072],
            prg05[3055:3040],prg05[3023:3008],prg05[2991:2976],prg05[2959:2944],prg05[2927:2912],prg05[2895:2880],prg05[2863:2848],prg05[2831:2816],
            prg05[2799:2784],prg05[2767:2752],prg05[2735:2720],prg05[2703:2688],prg05[2671:2656],prg05[2639:2624],prg05[2607:2592],prg05[2575:2560],
            prg05[2543:2528],prg05[2511:2496],prg05[2479:2464],prg05[2447:2432],prg05[2415:2400],prg05[2383:2368],prg05[2351:2336],prg05[2319:2304],
            prg05[2287:2272],prg05[2255:2240],prg05[2223:2208],prg05[2191:2176],prg05[2159:2144],prg05[2127:2112],prg05[2095:2080],prg05[2063:2048],
            prg05[2031:2016],prg05[1999:1984],prg05[1967:1952],prg05[1935:1920],prg05[1903:1888],prg05[1871:1856],prg05[1839:1824],prg05[1807:1792],
            prg05[1775:1760],prg05[1743:1728],prg05[1711:1696],prg05[1679:1664],prg05[1647:1632],prg05[1615:1600],prg05[1583:1568],prg05[1551:1536],
            prg05[1519:1504],prg05[1487:1472],prg05[1455:1440],prg05[1423:1408],prg05[1391:1376],prg05[1359:1344],prg05[1327:1312],prg05[1295:1280],
            prg05[1263:1248],prg05[1231:1216],prg05[1199:1184],prg05[1167:1152],prg05[1135:1120],prg05[1103:1088],prg05[1071:1056],prg05[1039:1024],
            prg05[1007: 992],prg05[ 975: 960],prg05[ 943: 928],prg05[ 911: 896],prg05[ 879: 864],prg05[ 847: 832],prg05[ 815: 800],prg05[ 783: 768],
            prg05[ 751: 736],prg05[ 719: 704],prg05[ 687: 672],prg05[ 655: 640],prg05[ 623: 608],prg05[ 591: 576],prg05[ 559: 544],prg05[ 527: 512],
            prg05[ 495: 480],prg05[ 463: 448],prg05[ 431: 416],prg05[ 399: 384],prg05[ 367: 352],prg05[ 335: 320],prg05[ 303: 288],prg05[ 271: 256],
            prg05[ 239: 224],prg05[ 207: 192],prg05[ 175: 160],prg05[ 143: 128],prg05[ 111:  96],prg05[  79:  64],prg05[  47:  32],prg05[  15:   0],
            prg04[4079:4064],prg04[4047:4032],prg04[4015:4000],prg04[3983:3968],prg04[3951:3936],prg04[3919:3904],prg04[3887:3872],prg04[3855:3840],
            prg04[3823:3808],prg04[3791:3776],prg04[3759:3744],prg04[3727:3712],prg04[3695:3680],prg04[3663:3648],prg04[3631:3616],prg04[3599:3584],
            prg04[3567:3552],prg04[3535:3520],prg04[3503:3488],prg04[3471:3456],prg04[3439:3424],prg04[3407:3392],prg04[3375:3360],prg04[3343:3328],
            prg04[3311:3296],prg04[3279:3264],prg04[3247:3232],prg04[3215:3200],prg04[3183:3168],prg04[3151:3136],prg04[3119:3104],prg04[3087:3072],
            prg04[3055:3040],prg04[3023:3008],prg04[2991:2976],prg04[2959:2944],prg04[2927:2912],prg04[2895:2880],prg04[2863:2848],prg04[2831:2816],
            prg04[2799:2784],prg04[2767:2752],prg04[2735:2720],prg04[2703:2688],prg04[2671:2656],prg04[2639:2624],prg04[2607:2592],prg04[2575:2560],
            prg04[2543:2528],prg04[2511:2496],prg04[2479:2464],prg04[2447:2432],prg04[2415:2400],prg04[2383:2368],prg04[2351:2336],prg04[2319:2304],
            prg04[2287:2272],prg04[2255:2240],prg04[2223:2208],prg04[2191:2176],prg04[2159:2144],prg04[2127:2112],prg04[2095:2080],prg04[2063:2048],
            prg04[2031:2016],prg04[1999:1984],prg04[1967:1952],prg04[1935:1920],prg04[1903:1888],prg04[1871:1856],prg04[1839:1824],prg04[1807:1792],
            prg04[1775:1760],prg04[1743:1728],prg04[1711:1696],prg04[1679:1664],prg04[1647:1632],prg04[1615:1600],prg04[1583:1568],prg04[1551:1536],
            prg04[1519:1504],prg04[1487:1472],prg04[1455:1440],prg04[1423:1408],prg04[1391:1376],prg04[1359:1344],prg04[1327:1312],prg04[1295:1280],
            prg04[1263:1248],prg04[1231:1216],prg04[1199:1184],prg04[1167:1152],prg04[1135:1120],prg04[1103:1088],prg04[1071:1056],prg04[1039:1024],
            prg04[1007: 992],prg04[ 975: 960],prg04[ 943: 928],prg04[ 911: 896],prg04[ 879: 864],prg04[ 847: 832],prg04[ 815: 800],prg04[ 783: 768],
            prg04[ 751: 736],prg04[ 719: 704],prg04[ 687: 672],prg04[ 655: 640],prg04[ 623: 608],prg04[ 591: 576],prg04[ 559: 544],prg04[ 527: 512],
            prg04[ 495: 480],prg04[ 463: 448],prg04[ 431: 416],prg04[ 399: 384],prg04[ 367: 352],prg04[ 335: 320],prg04[ 303: 288],prg04[ 271: 256],
            prg04[ 239: 224],prg04[ 207: 192],prg04[ 175: 160],prg04[ 143: 128],prg04[ 111:  96],prg04[  79:  64],prg04[  47:  32],prg04[  15:   0]};
   localparam [4095:0]
     pb1 = {prg03[4079:4064],prg03[4047:4032],prg03[4015:4000],prg03[3983:3968],prg03[3951:3936],prg03[3919:3904],prg03[3887:3872],prg03[3855:3840],
            prg03[3823:3808],prg03[3791:3776],prg03[3759:3744],prg03[3727:3712],prg03[3695:3680],prg03[3663:3648],prg03[3631:3616],prg03[3599:3584],
            prg03[3567:3552],prg03[3535:3520],prg03[3503:3488],prg03[3471:3456],prg03[3439:3424],prg03[3407:3392],prg03[3375:3360],prg03[3343:3328],
            prg03[3311:3296],prg03[3279:3264],prg03[3247:3232],prg03[3215:3200],prg03[3183:3168],prg03[3151:3136],prg03[3119:3104],prg03[3087:3072],
            prg03[3055:3040],prg03[3023:3008],prg03[2991:2976],prg03[2959:2944],prg03[2927:2912],prg03[2895:2880],prg03[2863:2848],prg03[2831:2816],
            prg03[2799:2784],prg03[2767:2752],prg03[2735:2720],prg03[2703:2688],prg03[2671:2656],prg03[2639:2624],prg03[2607:2592],prg03[2575:2560],
            prg03[2543:2528],prg03[2511:2496],prg03[2479:2464],prg03[2447:2432],prg03[2415:2400],prg03[2383:2368],prg03[2351:2336],prg03[2319:2304],
            prg03[2287:2272],prg03[2255:2240],prg03[2223:2208],prg03[2191:2176],prg03[2159:2144],prg03[2127:2112],prg03[2095:2080],prg03[2063:2048],
            prg03[2031:2016],prg03[1999:1984],prg03[1967:1952],prg03[1935:1920],prg03[1903:1888],prg03[1871:1856],prg03[1839:1824],prg03[1807:1792],
            prg03[1775:1760],prg03[1743:1728],prg03[1711:1696],prg03[1679:1664],prg03[1647:1632],prg03[1615:1600],prg03[1583:1568],prg03[1551:1536],
            prg03[1519:1504],prg03[1487:1472],prg03[1455:1440],prg03[1423:1408],prg03[1391:1376],prg03[1359:1344],prg03[1327:1312],prg03[1295:1280],
            prg03[1263:1248],prg03[1231:1216],prg03[1199:1184],prg03[1167:1152],prg03[1135:1120],prg03[1103:1088],prg03[1071:1056],prg03[1039:1024],
            prg03[1007: 992],prg03[ 975: 960],prg03[ 943: 928],prg03[ 911: 896],prg03[ 879: 864],prg03[ 847: 832],prg03[ 815: 800],prg03[ 783: 768],
            prg03[ 751: 736],prg03[ 719: 704],prg03[ 687: 672],prg03[ 655: 640],prg03[ 623: 608],prg03[ 591: 576],prg03[ 559: 544],prg03[ 527: 512],
            prg03[ 495: 480],prg03[ 463: 448],prg03[ 431: 416],prg03[ 399: 384],prg03[ 367: 352],prg03[ 335: 320],prg03[ 303: 288],prg03[ 271: 256],
            prg03[ 239: 224],prg03[ 207: 192],prg03[ 175: 160],prg03[ 143: 128],prg03[ 111:  96],prg03[  79:  64],prg03[  47:  32],prg03[  15:   0],
            prg02[4079:4064],prg02[4047:4032],prg02[4015:4000],prg02[3983:3968],prg02[3951:3936],prg02[3919:3904],prg02[3887:3872],prg02[3855:3840],
            prg02[3823:3808],prg02[3791:3776],prg02[3759:3744],prg02[3727:3712],prg02[3695:3680],prg02[3663:3648],prg02[3631:3616],prg02[3599:3584],
            prg02[3567:3552],prg02[3535:3520],prg02[3503:3488],prg02[3471:3456],prg02[3439:3424],prg02[3407:3392],prg02[3375:3360],prg02[3343:3328],
            prg02[3311:3296],prg02[3279:3264],prg02[3247:3232],prg02[3215:3200],prg02[3183:3168],prg02[3151:3136],prg02[3119:3104],prg02[3087:3072],
            prg02[3055:3040],prg02[3023:3008],prg02[2991:2976],prg02[2959:2944],prg02[2927:2912],prg02[2895:2880],prg02[2863:2848],prg02[2831:2816],
            prg02[2799:2784],prg02[2767:2752],prg02[2735:2720],prg02[2703:2688],prg02[2671:2656],prg02[2639:2624],prg02[2607:2592],prg02[2575:2560],
            prg02[2543:2528],prg02[2511:2496],prg02[2479:2464],prg02[2447:2432],prg02[2415:2400],prg02[2383:2368],prg02[2351:2336],prg02[2319:2304],
            prg02[2287:2272],prg02[2255:2240],prg02[2223:2208],prg02[2191:2176],prg02[2159:2144],prg02[2127:2112],prg02[2095:2080],prg02[2063:2048],
            prg02[2031:2016],prg02[1999:1984],prg02[1967:1952],prg02[1935:1920],prg02[1903:1888],prg02[1871:1856],prg02[1839:1824],prg02[1807:1792],
            prg02[1775:1760],prg02[1743:1728],prg02[1711:1696],prg02[1679:1664],prg02[1647:1632],prg02[1615:1600],prg02[1583:1568],prg02[1551:1536],
            prg02[1519:1504],prg02[1487:1472],prg02[1455:1440],prg02[1423:1408],prg02[1391:1376],prg02[1359:1344],prg02[1327:1312],prg02[1295:1280],
            prg02[1263:1248],prg02[1231:1216],prg02[1199:1184],prg02[1167:1152],prg02[1135:1120],prg02[1103:1088],prg02[1071:1056],prg02[1039:1024],
            prg02[1007: 992],prg02[ 975: 960],prg02[ 943: 928],prg02[ 911: 896],prg02[ 879: 864],prg02[ 847: 832],prg02[ 815: 800],prg02[ 783: 768],
            prg02[ 751: 736],prg02[ 719: 704],prg02[ 687: 672],prg02[ 655: 640],prg02[ 623: 608],prg02[ 591: 576],prg02[ 559: 544],prg02[ 527: 512],
            prg02[ 495: 480],prg02[ 463: 448],prg02[ 431: 416],prg02[ 399: 384],prg02[ 367: 352],prg02[ 335: 320],prg02[ 303: 288],prg02[ 271: 256],
            prg02[ 239: 224],prg02[ 207: 192],prg02[ 175: 160],prg02[ 143: 128],prg02[ 111:  96],prg02[  79:  64],prg02[  47:  32],prg02[  15:   0]};
   localparam [4095:0]
     pb0 = {prg01[4079:4064],prg01[4047:4032],prg01[4015:4000],prg01[3983:3968],prg01[3951:3936],prg01[3919:3904],prg01[3887:3872],prg01[3855:3840],
            prg01[3823:3808],prg01[3791:3776],prg01[3759:3744],prg01[3727:3712],prg01[3695:3680],prg01[3663:3648],prg01[3631:3616],prg01[3599:3584],
            prg01[3567:3552],prg01[3535:3520],prg01[3503:3488],prg01[3471:3456],prg01[3439:3424],prg01[3407:3392],prg01[3375:3360],prg01[3343:3328],
            prg01[3311:3296],prg01[3279:3264],prg01[3247:3232],prg01[3215:3200],prg01[3183:3168],prg01[3151:3136],prg01[3119:3104],prg01[3087:3072],
            prg01[3055:3040],prg01[3023:3008],prg01[2991:2976],prg01[2959:2944],prg01[2927:2912],prg01[2895:2880],prg01[2863:2848],prg01[2831:2816],
            prg01[2799:2784],prg01[2767:2752],prg01[2735:2720],prg01[2703:2688],prg01[2671:2656],prg01[2639:2624],prg01[2607:2592],prg01[2575:2560],
            prg01[2543:2528],prg01[2511:2496],prg01[2479:2464],prg01[2447:2432],prg01[2415:2400],prg01[2383:2368],prg01[2351:2336],prg01[2319:2304],
            prg01[2287:2272],prg01[2255:2240],prg01[2223:2208],prg01[2191:2176],prg01[2159:2144],prg01[2127:2112],prg01[2095:2080],prg01[2063:2048],
            prg01[2031:2016],prg01[1999:1984],prg01[1967:1952],prg01[1935:1920],prg01[1903:1888],prg01[1871:1856],prg01[1839:1824],prg01[1807:1792],
            prg01[1775:1760],prg01[1743:1728],prg01[1711:1696],prg01[1679:1664],prg01[1647:1632],prg01[1615:1600],prg01[1583:1568],prg01[1551:1536],
            prg01[1519:1504],prg01[1487:1472],prg01[1455:1440],prg01[1423:1408],prg01[1391:1376],prg01[1359:1344],prg01[1327:1312],prg01[1295:1280],
            prg01[1263:1248],prg01[1231:1216],prg01[1199:1184],prg01[1167:1152],prg01[1135:1120],prg01[1103:1088],prg01[1071:1056],prg01[1039:1024],
            prg01[1007: 992],prg01[ 975: 960],prg01[ 943: 928],prg01[ 911: 896],prg01[ 879: 864],prg01[ 847: 832],prg01[ 815: 800],prg01[ 783: 768],
            prg01[ 751: 736],prg01[ 719: 704],prg01[ 687: 672],prg01[ 655: 640],prg01[ 623: 608],prg01[ 591: 576],prg01[ 559: 544],prg01[ 527: 512],
            prg01[ 495: 480],prg01[ 463: 448],prg01[ 431: 416],prg01[ 399: 384],prg01[ 367: 352],prg01[ 335: 320],prg01[ 303: 288],prg01[ 271: 256],
            prg01[ 239: 224],prg01[ 207: 192],prg01[ 175: 160],prg01[ 143: 128],prg01[ 111:  96],prg01[  79:  64],prg01[  47:  32],prg01[  15:   0],
            prg00[4079:4064],prg00[4047:4032],prg00[4015:4000],prg00[3983:3968],prg00[3951:3936],prg00[3919:3904],prg00[3887:3872],prg00[3855:3840],
            prg00[3823:3808],prg00[3791:3776],prg00[3759:3744],prg00[3727:3712],prg00[3695:3680],prg00[3663:3648],prg00[3631:3616],prg00[3599:3584],
            prg00[3567:3552],prg00[3535:3520],prg00[3503:3488],prg00[3471:3456],prg00[3439:3424],prg00[3407:3392],prg00[3375:3360],prg00[3343:3328],
            prg00[3311:3296],prg00[3279:3264],prg00[3247:3232],prg00[3215:3200],prg00[3183:3168],prg00[3151:3136],prg00[3119:3104],prg00[3087:3072],
            prg00[3055:3040],prg00[3023:3008],prg00[2991:2976],prg00[2959:2944],prg00[2927:2912],prg00[2895:2880],prg00[2863:2848],prg00[2831:2816],
            prg00[2799:2784],prg00[2767:2752],prg00[2735:2720],prg00[2703:2688],prg00[2671:2656],prg00[2639:2624],prg00[2607:2592],prg00[2575:2560],
            prg00[2543:2528],prg00[2511:2496],prg00[2479:2464],prg00[2447:2432],prg00[2415:2400],prg00[2383:2368],prg00[2351:2336],prg00[2319:2304],
            prg00[2287:2272],prg00[2255:2240],prg00[2223:2208],prg00[2191:2176],prg00[2159:2144],prg00[2127:2112],prg00[2095:2080],prg00[2063:2048],
            prg00[2031:2016],prg00[1999:1984],prg00[1967:1952],prg00[1935:1920],prg00[1903:1888],prg00[1871:1856],prg00[1839:1824],prg00[1807:1792],
            prg00[1775:1760],prg00[1743:1728],prg00[1711:1696],prg00[1679:1664],prg00[1647:1632],prg00[1615:1600],prg00[1583:1568],prg00[1551:1536],
            prg00[1519:1504],prg00[1487:1472],prg00[1455:1440],prg00[1423:1408],prg00[1391:1376],prg00[1359:1344],prg00[1327:1312],prg00[1295:1280],
            prg00[1263:1248],prg00[1231:1216],prg00[1199:1184],prg00[1167:1152],prg00[1135:1120],prg00[1103:1088],prg00[1071:1056],prg00[1039:1024],
            prg00[1007: 992],prg00[ 975: 960],prg00[ 943: 928],prg00[ 911: 896],prg00[ 879: 864],prg00[ 847: 832],prg00[ 815: 800],prg00[ 783: 768],
            prg00[ 751: 736],prg00[ 719: 704],prg00[ 687: 672],prg00[ 655: 640],prg00[ 623: 608],prg00[ 591: 576],prg00[ 559: 544],prg00[ 527: 512],
            prg00[ 495: 480],prg00[ 463: 448],prg00[ 431: 416],prg00[ 399: 384],prg00[ 367: 352],prg00[ 335: 320],prg00[ 303: 288],prg00[ 271: 256],
            prg00[ 239: 224],prg00[ 207: 192],prg00[ 175: 160],prg00[ 143: 128],prg00[ 111:  96],prg00[  79:  64],prg00[  47:  32],prg00[  15:   0]};
   localparam [4095:0]
     ph7 = {prg0F[4095:4080],prg0F[4063:4048],prg0F[4031:4016],prg0F[3999:3984],prg0F[3967:3952],prg0F[3935:3920],prg0F[3903:3888],prg0F[3871:3856],
            prg0F[3839:3824],prg0F[3807:3792],prg0F[3775:3760],prg0F[3743:3728],prg0F[3711:3696],prg0F[3679:3664],prg0F[3647:3632],prg0F[3615:3600],
            prg0F[3583:3568],prg0F[3551:3536],prg0F[3519:3504],prg0F[3487:3472],prg0F[3455:3440],prg0F[3423:3408],prg0F[3391:3376],prg0F[3359:3344],
            prg0F[3327:3312],prg0F[3295:3280],prg0F[3263:3248],prg0F[3231:3216],prg0F[3199:3184],prg0F[3167:3152],prg0F[3135:3120],prg0F[3103:3088],
            prg0F[3071:3056],prg0F[3039:3024],prg0F[3007:2992],prg0F[2975:2960],prg0F[2943:2928],prg0F[2911:2896],prg0F[2879:2864],prg0F[2847:2832],
            prg0F[2815:2800],prg0F[2783:2768],prg0F[2751:2736],prg0F[2719:2704],prg0F[2687:2672],prg0F[2655:2640],prg0F[2623:2608],prg0F[2591:2576],
            prg0F[2559:2544],prg0F[2527:2512],prg0F[2495:2480],prg0F[2463:2448],prg0F[2431:2416],prg0F[2399:2384],prg0F[2367:2352],prg0F[2335:2320],
            prg0F[2303:2288],prg0F[2271:2256],prg0F[2239:2224],prg0F[2207:2192],prg0F[2175:2160],prg0F[2143:2128],prg0F[2111:2096],prg0F[2079:2064],
            prg0F[2047:2032],prg0F[2015:2000],prg0F[1983:1968],prg0F[1951:1936],prg0F[1919:1904],prg0F[1887:1872],prg0F[1855:1840],prg0F[1823:1808],
            prg0F[1791:1776],prg0F[1759:1744],prg0F[1727:1712],prg0F[1695:1680],prg0F[1663:1648],prg0F[1631:1616],prg0F[1599:1584],prg0F[1567:1552],
            prg0F[1535:1520],prg0F[1503:1488],prg0F[1471:1456],prg0F[1439:1424],prg0F[1407:1392],prg0F[1375:1360],prg0F[1343:1328],prg0F[1311:1296],
            prg0F[1279:1264],prg0F[1247:1232],prg0F[1215:1200],prg0F[1183:1168],prg0F[1151:1136],prg0F[1119:1104],prg0F[1087:1072],prg0F[1055:1040],
            prg0F[1023:1008],prg0F[ 991: 976],prg0F[ 959: 944],prg0F[ 927: 912],prg0F[ 895: 880],prg0F[ 863: 848],prg0F[ 831: 816],prg0F[ 799: 784],
            prg0F[ 767: 752],prg0F[ 735: 720],prg0F[ 703: 688],prg0F[ 671: 656],prg0F[ 639: 624],prg0F[ 607: 592],prg0F[ 575: 560],prg0F[ 543: 528],
            prg0F[ 511: 496],prg0F[ 479: 464],prg0F[ 447: 432],prg0F[ 415: 400],prg0F[ 383: 368],prg0F[ 351: 336],prg0F[ 319: 304],prg0F[ 287: 272],
            prg0F[ 255: 240],prg0F[ 223: 208],prg0F[ 191: 176],prg0F[ 159: 144],prg0F[ 127: 112],prg0F[  95:  80],prg0F[  63:  48],prg0F[  31:  16],
            prg0E[4095:4080],prg0E[4063:4048],prg0E[4031:4016],prg0E[3999:3984],prg0E[3967:3952],prg0E[3935:3920],prg0E[3903:3888],prg0E[3871:3856],
            prg0E[3839:3824],prg0E[3807:3792],prg0E[3775:3760],prg0E[3743:3728],prg0E[3711:3696],prg0E[3679:3664],prg0E[3647:3632],prg0E[3615:3600],
            prg0E[3583:3568],prg0E[3551:3536],prg0E[3519:3504],prg0E[3487:3472],prg0E[3455:3440],prg0E[3423:3408],prg0E[3391:3376],prg0E[3359:3344],
            prg0E[3327:3312],prg0E[3295:3280],prg0E[3263:3248],prg0E[3231:3216],prg0E[3199:3184],prg0E[3167:3152],prg0E[3135:3120],prg0E[3103:3088],
            prg0E[3071:3056],prg0E[3039:3024],prg0E[3007:2992],prg0E[2975:2960],prg0E[2943:2928],prg0E[2911:2896],prg0E[2879:2864],prg0E[2847:2832],
            prg0E[2815:2800],prg0E[2783:2768],prg0E[2751:2736],prg0E[2719:2704],prg0E[2687:2672],prg0E[2655:2640],prg0E[2623:2608],prg0E[2591:2576],
            prg0E[2559:2544],prg0E[2527:2512],prg0E[2495:2480],prg0E[2463:2448],prg0E[2431:2416],prg0E[2399:2384],prg0E[2367:2352],prg0E[2335:2320],
            prg0E[2303:2288],prg0E[2271:2256],prg0E[2239:2224],prg0E[2207:2192],prg0E[2175:2160],prg0E[2143:2128],prg0E[2111:2096],prg0E[2079:2064],
            prg0E[2047:2032],prg0E[2015:2000],prg0E[1983:1968],prg0E[1951:1936],prg0E[1919:1904],prg0E[1887:1872],prg0E[1855:1840],prg0E[1823:1808],
            prg0E[1791:1776],prg0E[1759:1744],prg0E[1727:1712],prg0E[1695:1680],prg0E[1663:1648],prg0E[1631:1616],prg0E[1599:1584],prg0E[1567:1552],
            prg0E[1535:1520],prg0E[1503:1488],prg0E[1471:1456],prg0E[1439:1424],prg0E[1407:1392],prg0E[1375:1360],prg0E[1343:1328],prg0E[1311:1296],
            prg0E[1279:1264],prg0E[1247:1232],prg0E[1215:1200],prg0E[1183:1168],prg0E[1151:1136],prg0E[1119:1104],prg0E[1087:1072],prg0E[1055:1040],
            prg0E[1023:1008],prg0E[ 991: 976],prg0E[ 959: 944],prg0E[ 927: 912],prg0E[ 895: 880],prg0E[ 863: 848],prg0E[ 831: 816],prg0E[ 799: 784],
            prg0E[ 767: 752],prg0E[ 735: 720],prg0E[ 703: 688],prg0E[ 671: 656],prg0E[ 639: 624],prg0E[ 607: 592],prg0E[ 575: 560],prg0E[ 543: 528],
            prg0E[ 511: 496],prg0E[ 479: 464],prg0E[ 447: 432],prg0E[ 415: 400],prg0E[ 383: 368],prg0E[ 351: 336],prg0E[ 319: 304],prg0E[ 287: 272],
            prg0E[ 255: 240],prg0E[ 223: 208],prg0E[ 191: 176],prg0E[ 159: 144],prg0E[ 127: 112],prg0E[  95:  80],prg0E[  63:  48],prg0E[  31:  16]};
   localparam [4095:0]
     ph6 = {prg0D[4095:4080],prg0D[4063:4048],prg0D[4031:4016],prg0D[3999:3984],prg0D[3967:3952],prg0D[3935:3920],prg0D[3903:3888],prg0D[3871:3856],
            prg0D[3839:3824],prg0D[3807:3792],prg0D[3775:3760],prg0D[3743:3728],prg0D[3711:3696],prg0D[3679:3664],prg0D[3647:3632],prg0D[3615:3600],
            prg0D[3583:3568],prg0D[3551:3536],prg0D[3519:3504],prg0D[3487:3472],prg0D[3455:3440],prg0D[3423:3408],prg0D[3391:3376],prg0D[3359:3344],
            prg0D[3327:3312],prg0D[3295:3280],prg0D[3263:3248],prg0D[3231:3216],prg0D[3199:3184],prg0D[3167:3152],prg0D[3135:3120],prg0D[3103:3088],
            prg0D[3071:3056],prg0D[3039:3024],prg0D[3007:2992],prg0D[2975:2960],prg0D[2943:2928],prg0D[2911:2896],prg0D[2879:2864],prg0D[2847:2832],
            prg0D[2815:2800],prg0D[2783:2768],prg0D[2751:2736],prg0D[2719:2704],prg0D[2687:2672],prg0D[2655:2640],prg0D[2623:2608],prg0D[2591:2576],
            prg0D[2559:2544],prg0D[2527:2512],prg0D[2495:2480],prg0D[2463:2448],prg0D[2431:2416],prg0D[2399:2384],prg0D[2367:2352],prg0D[2335:2320],
            prg0D[2303:2288],prg0D[2271:2256],prg0D[2239:2224],prg0D[2207:2192],prg0D[2175:2160],prg0D[2143:2128],prg0D[2111:2096],prg0D[2079:2064],
            prg0D[2047:2032],prg0D[2015:2000],prg0D[1983:1968],prg0D[1951:1936],prg0D[1919:1904],prg0D[1887:1872],prg0D[1855:1840],prg0D[1823:1808],
            prg0D[1791:1776],prg0D[1759:1744],prg0D[1727:1712],prg0D[1695:1680],prg0D[1663:1648],prg0D[1631:1616],prg0D[1599:1584],prg0D[1567:1552],
            prg0D[1535:1520],prg0D[1503:1488],prg0D[1471:1456],prg0D[1439:1424],prg0D[1407:1392],prg0D[1375:1360],prg0D[1343:1328],prg0D[1311:1296],
            prg0D[1279:1264],prg0D[1247:1232],prg0D[1215:1200],prg0D[1183:1168],prg0D[1151:1136],prg0D[1119:1104],prg0D[1087:1072],prg0D[1055:1040],
            prg0D[1023:1008],prg0D[ 991: 976],prg0D[ 959: 944],prg0D[ 927: 912],prg0D[ 895: 880],prg0D[ 863: 848],prg0D[ 831: 816],prg0D[ 799: 784],
            prg0D[ 767: 752],prg0D[ 735: 720],prg0D[ 703: 688],prg0D[ 671: 656],prg0D[ 639: 624],prg0D[ 607: 592],prg0D[ 575: 560],prg0D[ 543: 528],
            prg0D[ 511: 496],prg0D[ 479: 464],prg0D[ 447: 432],prg0D[ 415: 400],prg0D[ 383: 368],prg0D[ 351: 336],prg0D[ 319: 304],prg0D[ 287: 272],
            prg0D[ 255: 240],prg0D[ 223: 208],prg0D[ 191: 176],prg0D[ 159: 144],prg0D[ 127: 112],prg0D[  95:  80],prg0D[  63:  48],prg0D[  31:  16],
            prg0C[4095:4080],prg0C[4063:4048],prg0C[4031:4016],prg0C[3999:3984],prg0C[3967:3952],prg0C[3935:3920],prg0C[3903:3888],prg0C[3871:3856],
            prg0C[3839:3824],prg0C[3807:3792],prg0C[3775:3760],prg0C[3743:3728],prg0C[3711:3696],prg0C[3679:3664],prg0C[3647:3632],prg0C[3615:3600],
            prg0C[3583:3568],prg0C[3551:3536],prg0C[3519:3504],prg0C[3487:3472],prg0C[3455:3440],prg0C[3423:3408],prg0C[3391:3376],prg0C[3359:3344],
            prg0C[3327:3312],prg0C[3295:3280],prg0C[3263:3248],prg0C[3231:3216],prg0C[3199:3184],prg0C[3167:3152],prg0C[3135:3120],prg0C[3103:3088],
            prg0C[3071:3056],prg0C[3039:3024],prg0C[3007:2992],prg0C[2975:2960],prg0C[2943:2928],prg0C[2911:2896],prg0C[2879:2864],prg0C[2847:2832],
            prg0C[2815:2800],prg0C[2783:2768],prg0C[2751:2736],prg0C[2719:2704],prg0C[2687:2672],prg0C[2655:2640],prg0C[2623:2608],prg0C[2591:2576],
            prg0C[2559:2544],prg0C[2527:2512],prg0C[2495:2480],prg0C[2463:2448],prg0C[2431:2416],prg0C[2399:2384],prg0C[2367:2352],prg0C[2335:2320],
            prg0C[2303:2288],prg0C[2271:2256],prg0C[2239:2224],prg0C[2207:2192],prg0C[2175:2160],prg0C[2143:2128],prg0C[2111:2096],prg0C[2079:2064],
            prg0C[2047:2032],prg0C[2015:2000],prg0C[1983:1968],prg0C[1951:1936],prg0C[1919:1904],prg0C[1887:1872],prg0C[1855:1840],prg0C[1823:1808],
            prg0C[1791:1776],prg0C[1759:1744],prg0C[1727:1712],prg0C[1695:1680],prg0C[1663:1648],prg0C[1631:1616],prg0C[1599:1584],prg0C[1567:1552],
            prg0C[1535:1520],prg0C[1503:1488],prg0C[1471:1456],prg0C[1439:1424],prg0C[1407:1392],prg0C[1375:1360],prg0C[1343:1328],prg0C[1311:1296],
            prg0C[1279:1264],prg0C[1247:1232],prg0C[1215:1200],prg0C[1183:1168],prg0C[1151:1136],prg0C[1119:1104],prg0C[1087:1072],prg0C[1055:1040],
            prg0C[1023:1008],prg0C[ 991: 976],prg0C[ 959: 944],prg0C[ 927: 912],prg0C[ 895: 880],prg0C[ 863: 848],prg0C[ 831: 816],prg0C[ 799: 784],
            prg0C[ 767: 752],prg0C[ 735: 720],prg0C[ 703: 688],prg0C[ 671: 656],prg0C[ 639: 624],prg0C[ 607: 592],prg0C[ 575: 560],prg0C[ 543: 528],
            prg0C[ 511: 496],prg0C[ 479: 464],prg0C[ 447: 432],prg0C[ 415: 400],prg0C[ 383: 368],prg0C[ 351: 336],prg0C[ 319: 304],prg0C[ 287: 272],
            prg0C[ 255: 240],prg0C[ 223: 208],prg0C[ 191: 176],prg0C[ 159: 144],prg0C[ 127: 112],prg0C[  95:  80],prg0C[  63:  48],prg0C[  31:  16]};
   localparam [4095:0]
     ph5 = {prg0B[4095:4080],prg0B[4063:4048],prg0B[4031:4016],prg0B[3999:3984],prg0B[3967:3952],prg0B[3935:3920],prg0B[3903:3888],prg0B[3871:3856],
            prg0B[3839:3824],prg0B[3807:3792],prg0B[3775:3760],prg0B[3743:3728],prg0B[3711:3696],prg0B[3679:3664],prg0B[3647:3632],prg0B[3615:3600],
            prg0B[3583:3568],prg0B[3551:3536],prg0B[3519:3504],prg0B[3487:3472],prg0B[3455:3440],prg0B[3423:3408],prg0B[3391:3376],prg0B[3359:3344],
            prg0B[3327:3312],prg0B[3295:3280],prg0B[3263:3248],prg0B[3231:3216],prg0B[3199:3184],prg0B[3167:3152],prg0B[3135:3120],prg0B[3103:3088],
            prg0B[3071:3056],prg0B[3039:3024],prg0B[3007:2992],prg0B[2975:2960],prg0B[2943:2928],prg0B[2911:2896],prg0B[2879:2864],prg0B[2847:2832],
            prg0B[2815:2800],prg0B[2783:2768],prg0B[2751:2736],prg0B[2719:2704],prg0B[2687:2672],prg0B[2655:2640],prg0B[2623:2608],prg0B[2591:2576],
            prg0B[2559:2544],prg0B[2527:2512],prg0B[2495:2480],prg0B[2463:2448],prg0B[2431:2416],prg0B[2399:2384],prg0B[2367:2352],prg0B[2335:2320],
            prg0B[2303:2288],prg0B[2271:2256],prg0B[2239:2224],prg0B[2207:2192],prg0B[2175:2160],prg0B[2143:2128],prg0B[2111:2096],prg0B[2079:2064],
            prg0B[2047:2032],prg0B[2015:2000],prg0B[1983:1968],prg0B[1951:1936],prg0B[1919:1904],prg0B[1887:1872],prg0B[1855:1840],prg0B[1823:1808],
            prg0B[1791:1776],prg0B[1759:1744],prg0B[1727:1712],prg0B[1695:1680],prg0B[1663:1648],prg0B[1631:1616],prg0B[1599:1584],prg0B[1567:1552],
            prg0B[1535:1520],prg0B[1503:1488],prg0B[1471:1456],prg0B[1439:1424],prg0B[1407:1392],prg0B[1375:1360],prg0B[1343:1328],prg0B[1311:1296],
            prg0B[1279:1264],prg0B[1247:1232],prg0B[1215:1200],prg0B[1183:1168],prg0B[1151:1136],prg0B[1119:1104],prg0B[1087:1072],prg0B[1055:1040],
            prg0B[1023:1008],prg0B[ 991: 976],prg0B[ 959: 944],prg0B[ 927: 912],prg0B[ 895: 880],prg0B[ 863: 848],prg0B[ 831: 816],prg0B[ 799: 784],
            prg0B[ 767: 752],prg0B[ 735: 720],prg0B[ 703: 688],prg0B[ 671: 656],prg0B[ 639: 624],prg0B[ 607: 592],prg0B[ 575: 560],prg0B[ 543: 528],
            prg0B[ 511: 496],prg0B[ 479: 464],prg0B[ 447: 432],prg0B[ 415: 400],prg0B[ 383: 368],prg0B[ 351: 336],prg0B[ 319: 304],prg0B[ 287: 272],
            prg0B[ 255: 240],prg0B[ 223: 208],prg0B[ 191: 176],prg0B[ 159: 144],prg0B[ 127: 112],prg0B[  95:  80],prg0B[  63:  48],prg0B[  31:  16],
            prg0A[4095:4080],prg0A[4063:4048],prg0A[4031:4016],prg0A[3999:3984],prg0A[3967:3952],prg0A[3935:3920],prg0A[3903:3888],prg0A[3871:3856],
            prg0A[3839:3824],prg0A[3807:3792],prg0A[3775:3760],prg0A[3743:3728],prg0A[3711:3696],prg0A[3679:3664],prg0A[3647:3632],prg0A[3615:3600],
            prg0A[3583:3568],prg0A[3551:3536],prg0A[3519:3504],prg0A[3487:3472],prg0A[3455:3440],prg0A[3423:3408],prg0A[3391:3376],prg0A[3359:3344],
            prg0A[3327:3312],prg0A[3295:3280],prg0A[3263:3248],prg0A[3231:3216],prg0A[3199:3184],prg0A[3167:3152],prg0A[3135:3120],prg0A[3103:3088],
            prg0A[3071:3056],prg0A[3039:3024],prg0A[3007:2992],prg0A[2975:2960],prg0A[2943:2928],prg0A[2911:2896],prg0A[2879:2864],prg0A[2847:2832],
            prg0A[2815:2800],prg0A[2783:2768],prg0A[2751:2736],prg0A[2719:2704],prg0A[2687:2672],prg0A[2655:2640],prg0A[2623:2608],prg0A[2591:2576],
            prg0A[2559:2544],prg0A[2527:2512],prg0A[2495:2480],prg0A[2463:2448],prg0A[2431:2416],prg0A[2399:2384],prg0A[2367:2352],prg0A[2335:2320],
            prg0A[2303:2288],prg0A[2271:2256],prg0A[2239:2224],prg0A[2207:2192],prg0A[2175:2160],prg0A[2143:2128],prg0A[2111:2096],prg0A[2079:2064],
            prg0A[2047:2032],prg0A[2015:2000],prg0A[1983:1968],prg0A[1951:1936],prg0A[1919:1904],prg0A[1887:1872],prg0A[1855:1840],prg0A[1823:1808],
            prg0A[1791:1776],prg0A[1759:1744],prg0A[1727:1712],prg0A[1695:1680],prg0A[1663:1648],prg0A[1631:1616],prg0A[1599:1584],prg0A[1567:1552],
            prg0A[1535:1520],prg0A[1503:1488],prg0A[1471:1456],prg0A[1439:1424],prg0A[1407:1392],prg0A[1375:1360],prg0A[1343:1328],prg0A[1311:1296],
            prg0A[1279:1264],prg0A[1247:1232],prg0A[1215:1200],prg0A[1183:1168],prg0A[1151:1136],prg0A[1119:1104],prg0A[1087:1072],prg0A[1055:1040],
            prg0A[1023:1008],prg0A[ 991: 976],prg0A[ 959: 944],prg0A[ 927: 912],prg0A[ 895: 880],prg0A[ 863: 848],prg0A[ 831: 816],prg0A[ 799: 784],
            prg0A[ 767: 752],prg0A[ 735: 720],prg0A[ 703: 688],prg0A[ 671: 656],prg0A[ 639: 624],prg0A[ 607: 592],prg0A[ 575: 560],prg0A[ 543: 528],
            prg0A[ 511: 496],prg0A[ 479: 464],prg0A[ 447: 432],prg0A[ 415: 400],prg0A[ 383: 368],prg0A[ 351: 336],prg0A[ 319: 304],prg0A[ 287: 272],
            prg0A[ 255: 240],prg0A[ 223: 208],prg0A[ 191: 176],prg0A[ 159: 144],prg0A[ 127: 112],prg0A[  95:  80],prg0A[  63:  48],prg0A[  31:  16]};
   localparam [4095:0]
     ph4 = {prg09[4095:4080],prg09[4063:4048],prg09[4031:4016],prg09[3999:3984],prg09[3967:3952],prg09[3935:3920],prg09[3903:3888],prg09[3871:3856],
            prg09[3839:3824],prg09[3807:3792],prg09[3775:3760],prg09[3743:3728],prg09[3711:3696],prg09[3679:3664],prg09[3647:3632],prg09[3615:3600],
            prg09[3583:3568],prg09[3551:3536],prg09[3519:3504],prg09[3487:3472],prg09[3455:3440],prg09[3423:3408],prg09[3391:3376],prg09[3359:3344],
            prg09[3327:3312],prg09[3295:3280],prg09[3263:3248],prg09[3231:3216],prg09[3199:3184],prg09[3167:3152],prg09[3135:3120],prg09[3103:3088],
            prg09[3071:3056],prg09[3039:3024],prg09[3007:2992],prg09[2975:2960],prg09[2943:2928],prg09[2911:2896],prg09[2879:2864],prg09[2847:2832],
            prg09[2815:2800],prg09[2783:2768],prg09[2751:2736],prg09[2719:2704],prg09[2687:2672],prg09[2655:2640],prg09[2623:2608],prg09[2591:2576],
            prg09[2559:2544],prg09[2527:2512],prg09[2495:2480],prg09[2463:2448],prg09[2431:2416],prg09[2399:2384],prg09[2367:2352],prg09[2335:2320],
            prg09[2303:2288],prg09[2271:2256],prg09[2239:2224],prg09[2207:2192],prg09[2175:2160],prg09[2143:2128],prg09[2111:2096],prg09[2079:2064],
            prg09[2047:2032],prg09[2015:2000],prg09[1983:1968],prg09[1951:1936],prg09[1919:1904],prg09[1887:1872],prg09[1855:1840],prg09[1823:1808],
            prg09[1791:1776],prg09[1759:1744],prg09[1727:1712],prg09[1695:1680],prg09[1663:1648],prg09[1631:1616],prg09[1599:1584],prg09[1567:1552],
            prg09[1535:1520],prg09[1503:1488],prg09[1471:1456],prg09[1439:1424],prg09[1407:1392],prg09[1375:1360],prg09[1343:1328],prg09[1311:1296],
            prg09[1279:1264],prg09[1247:1232],prg09[1215:1200],prg09[1183:1168],prg09[1151:1136],prg09[1119:1104],prg09[1087:1072],prg09[1055:1040],
            prg09[1023:1008],prg09[ 991: 976],prg09[ 959: 944],prg09[ 927: 912],prg09[ 895: 880],prg09[ 863: 848],prg09[ 831: 816],prg09[ 799: 784],
            prg09[ 767: 752],prg09[ 735: 720],prg09[ 703: 688],prg09[ 671: 656],prg09[ 639: 624],prg09[ 607: 592],prg09[ 575: 560],prg09[ 543: 528],
            prg09[ 511: 496],prg09[ 479: 464],prg09[ 447: 432],prg09[ 415: 400],prg09[ 383: 368],prg09[ 351: 336],prg09[ 319: 304],prg09[ 287: 272],
            prg09[ 255: 240],prg09[ 223: 208],prg09[ 191: 176],prg09[ 159: 144],prg09[ 127: 112],prg09[  95:  80],prg09[  63:  48],prg09[  31:  16],
            prg08[4095:4080],prg08[4063:4048],prg08[4031:4016],prg08[3999:3984],prg08[3967:3952],prg08[3935:3920],prg08[3903:3888],prg08[3871:3856],
            prg08[3839:3824],prg08[3807:3792],prg08[3775:3760],prg08[3743:3728],prg08[3711:3696],prg08[3679:3664],prg08[3647:3632],prg08[3615:3600],
            prg08[3583:3568],prg08[3551:3536],prg08[3519:3504],prg08[3487:3472],prg08[3455:3440],prg08[3423:3408],prg08[3391:3376],prg08[3359:3344],
            prg08[3327:3312],prg08[3295:3280],prg08[3263:3248],prg08[3231:3216],prg08[3199:3184],prg08[3167:3152],prg08[3135:3120],prg08[3103:3088],
            prg08[3071:3056],prg08[3039:3024],prg08[3007:2992],prg08[2975:2960],prg08[2943:2928],prg08[2911:2896],prg08[2879:2864],prg08[2847:2832],
            prg08[2815:2800],prg08[2783:2768],prg08[2751:2736],prg08[2719:2704],prg08[2687:2672],prg08[2655:2640],prg08[2623:2608],prg08[2591:2576],
            prg08[2559:2544],prg08[2527:2512],prg08[2495:2480],prg08[2463:2448],prg08[2431:2416],prg08[2399:2384],prg08[2367:2352],prg08[2335:2320],
            prg08[2303:2288],prg08[2271:2256],prg08[2239:2224],prg08[2207:2192],prg08[2175:2160],prg08[2143:2128],prg08[2111:2096],prg08[2079:2064],
            prg08[2047:2032],prg08[2015:2000],prg08[1983:1968],prg08[1951:1936],prg08[1919:1904],prg08[1887:1872],prg08[1855:1840],prg08[1823:1808],
            prg08[1791:1776],prg08[1759:1744],prg08[1727:1712],prg08[1695:1680],prg08[1663:1648],prg08[1631:1616],prg08[1599:1584],prg08[1567:1552],
            prg08[1535:1520],prg08[1503:1488],prg08[1471:1456],prg08[1439:1424],prg08[1407:1392],prg08[1375:1360],prg08[1343:1328],prg08[1311:1296],
            prg08[1279:1264],prg08[1247:1232],prg08[1215:1200],prg08[1183:1168],prg08[1151:1136],prg08[1119:1104],prg08[1087:1072],prg08[1055:1040],
            prg08[1023:1008],prg08[ 991: 976],prg08[ 959: 944],prg08[ 927: 912],prg08[ 895: 880],prg08[ 863: 848],prg08[ 831: 816],prg08[ 799: 784],
            prg08[ 767: 752],prg08[ 735: 720],prg08[ 703: 688],prg08[ 671: 656],prg08[ 639: 624],prg08[ 607: 592],prg08[ 575: 560],prg08[ 543: 528],
            prg08[ 511: 496],prg08[ 479: 464],prg08[ 447: 432],prg08[ 415: 400],prg08[ 383: 368],prg08[ 351: 336],prg08[ 319: 304],prg08[ 287: 272],
            prg08[ 255: 240],prg08[ 223: 208],prg08[ 191: 176],prg08[ 159: 144],prg08[ 127: 112],prg08[  95:  80],prg08[  63:  48],prg08[  31:  16]};
   localparam [4095:0]
     ph3 = {prg07[4095:4080],prg07[4063:4048],prg07[4031:4016],prg07[3999:3984],prg07[3967:3952],prg07[3935:3920],prg07[3903:3888],prg07[3871:3856],
            prg07[3839:3824],prg07[3807:3792],prg07[3775:3760],prg07[3743:3728],prg07[3711:3696],prg07[3679:3664],prg07[3647:3632],prg07[3615:3600],
            prg07[3583:3568],prg07[3551:3536],prg07[3519:3504],prg07[3487:3472],prg07[3455:3440],prg07[3423:3408],prg07[3391:3376],prg07[3359:3344],
            prg07[3327:3312],prg07[3295:3280],prg07[3263:3248],prg07[3231:3216],prg07[3199:3184],prg07[3167:3152],prg07[3135:3120],prg07[3103:3088],
            prg07[3071:3056],prg07[3039:3024],prg07[3007:2992],prg07[2975:2960],prg07[2943:2928],prg07[2911:2896],prg07[2879:2864],prg07[2847:2832],
            prg07[2815:2800],prg07[2783:2768],prg07[2751:2736],prg07[2719:2704],prg07[2687:2672],prg07[2655:2640],prg07[2623:2608],prg07[2591:2576],
            prg07[2559:2544],prg07[2527:2512],prg07[2495:2480],prg07[2463:2448],prg07[2431:2416],prg07[2399:2384],prg07[2367:2352],prg07[2335:2320],
            prg07[2303:2288],prg07[2271:2256],prg07[2239:2224],prg07[2207:2192],prg07[2175:2160],prg07[2143:2128],prg07[2111:2096],prg07[2079:2064],
            prg07[2047:2032],prg07[2015:2000],prg07[1983:1968],prg07[1951:1936],prg07[1919:1904],prg07[1887:1872],prg07[1855:1840],prg07[1823:1808],
            prg07[1791:1776],prg07[1759:1744],prg07[1727:1712],prg07[1695:1680],prg07[1663:1648],prg07[1631:1616],prg07[1599:1584],prg07[1567:1552],
            prg07[1535:1520],prg07[1503:1488],prg07[1471:1456],prg07[1439:1424],prg07[1407:1392],prg07[1375:1360],prg07[1343:1328],prg07[1311:1296],
            prg07[1279:1264],prg07[1247:1232],prg07[1215:1200],prg07[1183:1168],prg07[1151:1136],prg07[1119:1104],prg07[1087:1072],prg07[1055:1040],
            prg07[1023:1008],prg07[ 991: 976],prg07[ 959: 944],prg07[ 927: 912],prg07[ 895: 880],prg07[ 863: 848],prg07[ 831: 816],prg07[ 799: 784],
            prg07[ 767: 752],prg07[ 735: 720],prg07[ 703: 688],prg07[ 671: 656],prg07[ 639: 624],prg07[ 607: 592],prg07[ 575: 560],prg07[ 543: 528],
            prg07[ 511: 496],prg07[ 479: 464],prg07[ 447: 432],prg07[ 415: 400],prg07[ 383: 368],prg07[ 351: 336],prg07[ 319: 304],prg07[ 287: 272],
            prg07[ 255: 240],prg07[ 223: 208],prg07[ 191: 176],prg07[ 159: 144],prg07[ 127: 112],prg07[  95:  80],prg07[  63:  48],prg07[  31:  16],
            prg06[4095:4080],prg06[4063:4048],prg06[4031:4016],prg06[3999:3984],prg06[3967:3952],prg06[3935:3920],prg06[3903:3888],prg06[3871:3856],
            prg06[3839:3824],prg06[3807:3792],prg06[3775:3760],prg06[3743:3728],prg06[3711:3696],prg06[3679:3664],prg06[3647:3632],prg06[3615:3600],
            prg06[3583:3568],prg06[3551:3536],prg06[3519:3504],prg06[3487:3472],prg06[3455:3440],prg06[3423:3408],prg06[3391:3376],prg06[3359:3344],
            prg06[3327:3312],prg06[3295:3280],prg06[3263:3248],prg06[3231:3216],prg06[3199:3184],prg06[3167:3152],prg06[3135:3120],prg06[3103:3088],
            prg06[3071:3056],prg06[3039:3024],prg06[3007:2992],prg06[2975:2960],prg06[2943:2928],prg06[2911:2896],prg06[2879:2864],prg06[2847:2832],
            prg06[2815:2800],prg06[2783:2768],prg06[2751:2736],prg06[2719:2704],prg06[2687:2672],prg06[2655:2640],prg06[2623:2608],prg06[2591:2576],
            prg06[2559:2544],prg06[2527:2512],prg06[2495:2480],prg06[2463:2448],prg06[2431:2416],prg06[2399:2384],prg06[2367:2352],prg06[2335:2320],
            prg06[2303:2288],prg06[2271:2256],prg06[2239:2224],prg06[2207:2192],prg06[2175:2160],prg06[2143:2128],prg06[2111:2096],prg06[2079:2064],
            prg06[2047:2032],prg06[2015:2000],prg06[1983:1968],prg06[1951:1936],prg06[1919:1904],prg06[1887:1872],prg06[1855:1840],prg06[1823:1808],
            prg06[1791:1776],prg06[1759:1744],prg06[1727:1712],prg06[1695:1680],prg06[1663:1648],prg06[1631:1616],prg06[1599:1584],prg06[1567:1552],
            prg06[1535:1520],prg06[1503:1488],prg06[1471:1456],prg06[1439:1424],prg06[1407:1392],prg06[1375:1360],prg06[1343:1328],prg06[1311:1296],
            prg06[1279:1264],prg06[1247:1232],prg06[1215:1200],prg06[1183:1168],prg06[1151:1136],prg06[1119:1104],prg06[1087:1072],prg06[1055:1040],
            prg06[1023:1008],prg06[ 991: 976],prg06[ 959: 944],prg06[ 927: 912],prg06[ 895: 880],prg06[ 863: 848],prg06[ 831: 816],prg06[ 799: 784],
            prg06[ 767: 752],prg06[ 735: 720],prg06[ 703: 688],prg06[ 671: 656],prg06[ 639: 624],prg06[ 607: 592],prg06[ 575: 560],prg06[ 543: 528],
            prg06[ 511: 496],prg06[ 479: 464],prg06[ 447: 432],prg06[ 415: 400],prg06[ 383: 368],prg06[ 351: 336],prg06[ 319: 304],prg06[ 287: 272],
            prg06[ 255: 240],prg06[ 223: 208],prg06[ 191: 176],prg06[ 159: 144],prg06[ 127: 112],prg06[  95:  80],prg06[  63:  48],prg06[  31:  16]};
   localparam [4095:0]
     ph2 = {prg05[4095:4080],prg05[4063:4048],prg05[4031:4016],prg05[3999:3984],prg05[3967:3952],prg05[3935:3920],prg05[3903:3888],prg05[3871:3856],
            prg05[3839:3824],prg05[3807:3792],prg05[3775:3760],prg05[3743:3728],prg05[3711:3696],prg05[3679:3664],prg05[3647:3632],prg05[3615:3600],
            prg05[3583:3568],prg05[3551:3536],prg05[3519:3504],prg05[3487:3472],prg05[3455:3440],prg05[3423:3408],prg05[3391:3376],prg05[3359:3344],
            prg05[3327:3312],prg05[3295:3280],prg05[3263:3248],prg05[3231:3216],prg05[3199:3184],prg05[3167:3152],prg05[3135:3120],prg05[3103:3088],
            prg05[3071:3056],prg05[3039:3024],prg05[3007:2992],prg05[2975:2960],prg05[2943:2928],prg05[2911:2896],prg05[2879:2864],prg05[2847:2832],
            prg05[2815:2800],prg05[2783:2768],prg05[2751:2736],prg05[2719:2704],prg05[2687:2672],prg05[2655:2640],prg05[2623:2608],prg05[2591:2576],
            prg05[2559:2544],prg05[2527:2512],prg05[2495:2480],prg05[2463:2448],prg05[2431:2416],prg05[2399:2384],prg05[2367:2352],prg05[2335:2320],
            prg05[2303:2288],prg05[2271:2256],prg05[2239:2224],prg05[2207:2192],prg05[2175:2160],prg05[2143:2128],prg05[2111:2096],prg05[2079:2064],
            prg05[2047:2032],prg05[2015:2000],prg05[1983:1968],prg05[1951:1936],prg05[1919:1904],prg05[1887:1872],prg05[1855:1840],prg05[1823:1808],
            prg05[1791:1776],prg05[1759:1744],prg05[1727:1712],prg05[1695:1680],prg05[1663:1648],prg05[1631:1616],prg05[1599:1584],prg05[1567:1552],
            prg05[1535:1520],prg05[1503:1488],prg05[1471:1456],prg05[1439:1424],prg05[1407:1392],prg05[1375:1360],prg05[1343:1328],prg05[1311:1296],
            prg05[1279:1264],prg05[1247:1232],prg05[1215:1200],prg05[1183:1168],prg05[1151:1136],prg05[1119:1104],prg05[1087:1072],prg05[1055:1040],
            prg05[1023:1008],prg05[ 991: 976],prg05[ 959: 944],prg05[ 927: 912],prg05[ 895: 880],prg05[ 863: 848],prg05[ 831: 816],prg05[ 799: 784],
            prg05[ 767: 752],prg05[ 735: 720],prg05[ 703: 688],prg05[ 671: 656],prg05[ 639: 624],prg05[ 607: 592],prg05[ 575: 560],prg05[ 543: 528],
            prg05[ 511: 496],prg05[ 479: 464],prg05[ 447: 432],prg05[ 415: 400],prg05[ 383: 368],prg05[ 351: 336],prg05[ 319: 304],prg05[ 287: 272],
            prg05[ 255: 240],prg05[ 223: 208],prg05[ 191: 176],prg05[ 159: 144],prg05[ 127: 112],prg05[  95:  80],prg05[  63:  48],prg05[  31:  16],
            prg04[4095:4080],prg04[4063:4048],prg04[4031:4016],prg04[3999:3984],prg04[3967:3952],prg04[3935:3920],prg04[3903:3888],prg04[3871:3856],
            prg04[3839:3824],prg04[3807:3792],prg04[3775:3760],prg04[3743:3728],prg04[3711:3696],prg04[3679:3664],prg04[3647:3632],prg04[3615:3600],
            prg04[3583:3568],prg04[3551:3536],prg04[3519:3504],prg04[3487:3472],prg04[3455:3440],prg04[3423:3408],prg04[3391:3376],prg04[3359:3344],
            prg04[3327:3312],prg04[3295:3280],prg04[3263:3248],prg04[3231:3216],prg04[3199:3184],prg04[3167:3152],prg04[3135:3120],prg04[3103:3088],
            prg04[3071:3056],prg04[3039:3024],prg04[3007:2992],prg04[2975:2960],prg04[2943:2928],prg04[2911:2896],prg04[2879:2864],prg04[2847:2832],
            prg04[2815:2800],prg04[2783:2768],prg04[2751:2736],prg04[2719:2704],prg04[2687:2672],prg04[2655:2640],prg04[2623:2608],prg04[2591:2576],
            prg04[2559:2544],prg04[2527:2512],prg04[2495:2480],prg04[2463:2448],prg04[2431:2416],prg04[2399:2384],prg04[2367:2352],prg04[2335:2320],
            prg04[2303:2288],prg04[2271:2256],prg04[2239:2224],prg04[2207:2192],prg04[2175:2160],prg04[2143:2128],prg04[2111:2096],prg04[2079:2064],
            prg04[2047:2032],prg04[2015:2000],prg04[1983:1968],prg04[1951:1936],prg04[1919:1904],prg04[1887:1872],prg04[1855:1840],prg04[1823:1808],
            prg04[1791:1776],prg04[1759:1744],prg04[1727:1712],prg04[1695:1680],prg04[1663:1648],prg04[1631:1616],prg04[1599:1584],prg04[1567:1552],
            prg04[1535:1520],prg04[1503:1488],prg04[1471:1456],prg04[1439:1424],prg04[1407:1392],prg04[1375:1360],prg04[1343:1328],prg04[1311:1296],
            prg04[1279:1264],prg04[1247:1232],prg04[1215:1200],prg04[1183:1168],prg04[1151:1136],prg04[1119:1104],prg04[1087:1072],prg04[1055:1040],
            prg04[1023:1008],prg04[ 991: 976],prg04[ 959: 944],prg04[ 927: 912],prg04[ 895: 880],prg04[ 863: 848],prg04[ 831: 816],prg04[ 799: 784],
            prg04[ 767: 752],prg04[ 735: 720],prg04[ 703: 688],prg04[ 671: 656],prg04[ 639: 624],prg04[ 607: 592],prg04[ 575: 560],prg04[ 543: 528],
            prg04[ 511: 496],prg04[ 479: 464],prg04[ 447: 432],prg04[ 415: 400],prg04[ 383: 368],prg04[ 351: 336],prg04[ 319: 304],prg04[ 287: 272],
            prg04[ 255: 240],prg04[ 223: 208],prg04[ 191: 176],prg04[ 159: 144],prg04[ 127: 112],prg04[  95:  80],prg04[  63:  48],prg04[  31:  16]};
   localparam [4095:0]
     ph1 = {prg03[4095:4080],prg03[4063:4048],prg03[4031:4016],prg03[3999:3984],prg03[3967:3952],prg03[3935:3920],prg03[3903:3888],prg03[3871:3856],
            prg03[3839:3824],prg03[3807:3792],prg03[3775:3760],prg03[3743:3728],prg03[3711:3696],prg03[3679:3664],prg03[3647:3632],prg03[3615:3600],
            prg03[3583:3568],prg03[3551:3536],prg03[3519:3504],prg03[3487:3472],prg03[3455:3440],prg03[3423:3408],prg03[3391:3376],prg03[3359:3344],
            prg03[3327:3312],prg03[3295:3280],prg03[3263:3248],prg03[3231:3216],prg03[3199:3184],prg03[3167:3152],prg03[3135:3120],prg03[3103:3088],
            prg03[3071:3056],prg03[3039:3024],prg03[3007:2992],prg03[2975:2960],prg03[2943:2928],prg03[2911:2896],prg03[2879:2864],prg03[2847:2832],
            prg03[2815:2800],prg03[2783:2768],prg03[2751:2736],prg03[2719:2704],prg03[2687:2672],prg03[2655:2640],prg03[2623:2608],prg03[2591:2576],
            prg03[2559:2544],prg03[2527:2512],prg03[2495:2480],prg03[2463:2448],prg03[2431:2416],prg03[2399:2384],prg03[2367:2352],prg03[2335:2320],
            prg03[2303:2288],prg03[2271:2256],prg03[2239:2224],prg03[2207:2192],prg03[2175:2160],prg03[2143:2128],prg03[2111:2096],prg03[2079:2064],
            prg03[2047:2032],prg03[2015:2000],prg03[1983:1968],prg03[1951:1936],prg03[1919:1904],prg03[1887:1872],prg03[1855:1840],prg03[1823:1808],
            prg03[1791:1776],prg03[1759:1744],prg03[1727:1712],prg03[1695:1680],prg03[1663:1648],prg03[1631:1616],prg03[1599:1584],prg03[1567:1552],
            prg03[1535:1520],prg03[1503:1488],prg03[1471:1456],prg03[1439:1424],prg03[1407:1392],prg03[1375:1360],prg03[1343:1328],prg03[1311:1296],
            prg03[1279:1264],prg03[1247:1232],prg03[1215:1200],prg03[1183:1168],prg03[1151:1136],prg03[1119:1104],prg03[1087:1072],prg03[1055:1040],
            prg03[1023:1008],prg03[ 991: 976],prg03[ 959: 944],prg03[ 927: 912],prg03[ 895: 880],prg03[ 863: 848],prg03[ 831: 816],prg03[ 799: 784],
            prg03[ 767: 752],prg03[ 735: 720],prg03[ 703: 688],prg03[ 671: 656],prg03[ 639: 624],prg03[ 607: 592],prg03[ 575: 560],prg03[ 543: 528],
            prg03[ 511: 496],prg03[ 479: 464],prg03[ 447: 432],prg03[ 415: 400],prg03[ 383: 368],prg03[ 351: 336],prg03[ 319: 304],prg03[ 287: 272],
            prg03[ 255: 240],prg03[ 223: 208],prg03[ 191: 176],prg03[ 159: 144],prg03[ 127: 112],prg03[  95:  80],prg03[  63:  48],prg03[  31:  16],
            prg02[4095:4080],prg02[4063:4048],prg02[4031:4016],prg02[3999:3984],prg02[3967:3952],prg02[3935:3920],prg02[3903:3888],prg02[3871:3856],
            prg02[3839:3824],prg02[3807:3792],prg02[3775:3760],prg02[3743:3728],prg02[3711:3696],prg02[3679:3664],prg02[3647:3632],prg02[3615:3600],
            prg02[3583:3568],prg02[3551:3536],prg02[3519:3504],prg02[3487:3472],prg02[3455:3440],prg02[3423:3408],prg02[3391:3376],prg02[3359:3344],
            prg02[3327:3312],prg02[3295:3280],prg02[3263:3248],prg02[3231:3216],prg02[3199:3184],prg02[3167:3152],prg02[3135:3120],prg02[3103:3088],
            prg02[3071:3056],prg02[3039:3024],prg02[3007:2992],prg02[2975:2960],prg02[2943:2928],prg02[2911:2896],prg02[2879:2864],prg02[2847:2832],
            prg02[2815:2800],prg02[2783:2768],prg02[2751:2736],prg02[2719:2704],prg02[2687:2672],prg02[2655:2640],prg02[2623:2608],prg02[2591:2576],
            prg02[2559:2544],prg02[2527:2512],prg02[2495:2480],prg02[2463:2448],prg02[2431:2416],prg02[2399:2384],prg02[2367:2352],prg02[2335:2320],
            prg02[2303:2288],prg02[2271:2256],prg02[2239:2224],prg02[2207:2192],prg02[2175:2160],prg02[2143:2128],prg02[2111:2096],prg02[2079:2064],
            prg02[2047:2032],prg02[2015:2000],prg02[1983:1968],prg02[1951:1936],prg02[1919:1904],prg02[1887:1872],prg02[1855:1840],prg02[1823:1808],
            prg02[1791:1776],prg02[1759:1744],prg02[1727:1712],prg02[1695:1680],prg02[1663:1648],prg02[1631:1616],prg02[1599:1584],prg02[1567:1552],
            prg02[1535:1520],prg02[1503:1488],prg02[1471:1456],prg02[1439:1424],prg02[1407:1392],prg02[1375:1360],prg02[1343:1328],prg02[1311:1296],
            prg02[1279:1264],prg02[1247:1232],prg02[1215:1200],prg02[1183:1168],prg02[1151:1136],prg02[1119:1104],prg02[1087:1072],prg02[1055:1040],
            prg02[1023:1008],prg02[ 991: 976],prg02[ 959: 944],prg02[ 927: 912],prg02[ 895: 880],prg02[ 863: 848],prg02[ 831: 816],prg02[ 799: 784],
            prg02[ 767: 752],prg02[ 735: 720],prg02[ 703: 688],prg02[ 671: 656],prg02[ 639: 624],prg02[ 607: 592],prg02[ 575: 560],prg02[ 543: 528],
            prg02[ 511: 496],prg02[ 479: 464],prg02[ 447: 432],prg02[ 415: 400],prg02[ 383: 368],prg02[ 351: 336],prg02[ 319: 304],prg02[ 287: 272],
            prg02[ 255: 240],prg02[ 223: 208],prg02[ 191: 176],prg02[ 159: 144],prg02[ 127: 112],prg02[  95:  80],prg02[  63:  48],prg02[  31:  16]};
   localparam [4095:0]
     ph0 = {prg01[4095:4080],prg01[4063:4048],prg01[4031:4016],prg01[3999:3984],prg01[3967:3952],prg01[3935:3920],prg01[3903:3888],prg01[3871:3856],
            prg01[3839:3824],prg01[3807:3792],prg01[3775:3760],prg01[3743:3728],prg01[3711:3696],prg01[3679:3664],prg01[3647:3632],prg01[3615:3600],
            prg01[3583:3568],prg01[3551:3536],prg01[3519:3504],prg01[3487:3472],prg01[3455:3440],prg01[3423:3408],prg01[3391:3376],prg01[3359:3344],
            prg01[3327:3312],prg01[3295:3280],prg01[3263:3248],prg01[3231:3216],prg01[3199:3184],prg01[3167:3152],prg01[3135:3120],prg01[3103:3088],
            prg01[3071:3056],prg01[3039:3024],prg01[3007:2992],prg01[2975:2960],prg01[2943:2928],prg01[2911:2896],prg01[2879:2864],prg01[2847:2832],
            prg01[2815:2800],prg01[2783:2768],prg01[2751:2736],prg01[2719:2704],prg01[2687:2672],prg01[2655:2640],prg01[2623:2608],prg01[2591:2576],
            prg01[2559:2544],prg01[2527:2512],prg01[2495:2480],prg01[2463:2448],prg01[2431:2416],prg01[2399:2384],prg01[2367:2352],prg01[2335:2320],
            prg01[2303:2288],prg01[2271:2256],prg01[2239:2224],prg01[2207:2192],prg01[2175:2160],prg01[2143:2128],prg01[2111:2096],prg01[2079:2064],
            prg01[2047:2032],prg01[2015:2000],prg01[1983:1968],prg01[1951:1936],prg01[1919:1904],prg01[1887:1872],prg01[1855:1840],prg01[1823:1808],
            prg01[1791:1776],prg01[1759:1744],prg01[1727:1712],prg01[1695:1680],prg01[1663:1648],prg01[1631:1616],prg01[1599:1584],prg01[1567:1552],
            prg01[1535:1520],prg01[1503:1488],prg01[1471:1456],prg01[1439:1424],prg01[1407:1392],prg01[1375:1360],prg01[1343:1328],prg01[1311:1296],
            prg01[1279:1264],prg01[1247:1232],prg01[1215:1200],prg01[1183:1168],prg01[1151:1136],prg01[1119:1104],prg01[1087:1072],prg01[1055:1040],
            prg01[1023:1008],prg01[ 991: 976],prg01[ 959: 944],prg01[ 927: 912],prg01[ 895: 880],prg01[ 863: 848],prg01[ 831: 816],prg01[ 799: 784],
            prg01[ 767: 752],prg01[ 735: 720],prg01[ 703: 688],prg01[ 671: 656],prg01[ 639: 624],prg01[ 607: 592],prg01[ 575: 560],prg01[ 543: 528],
            prg01[ 511: 496],prg01[ 479: 464],prg01[ 447: 432],prg01[ 415: 400],prg01[ 383: 368],prg01[ 351: 336],prg01[ 319: 304],prg01[ 287: 272],
            prg01[ 255: 240],prg01[ 223: 208],prg01[ 191: 176],prg01[ 159: 144],prg01[ 127: 112],prg01[  95:  80],prg01[  63:  48],prg01[  31:  16],
            prg00[4095:4080],prg00[4063:4048],prg00[4031:4016],prg00[3999:3984],prg00[3967:3952],prg00[3935:3920],prg00[3903:3888],prg00[3871:3856],
            prg00[3839:3824],prg00[3807:3792],prg00[3775:3760],prg00[3743:3728],prg00[3711:3696],prg00[3679:3664],prg00[3647:3632],prg00[3615:3600],
            prg00[3583:3568],prg00[3551:3536],prg00[3519:3504],prg00[3487:3472],prg00[3455:3440],prg00[3423:3408],prg00[3391:3376],prg00[3359:3344],
            prg00[3327:3312],prg00[3295:3280],prg00[3263:3248],prg00[3231:3216],prg00[3199:3184],prg00[3167:3152],prg00[3135:3120],prg00[3103:3088],
            prg00[3071:3056],prg00[3039:3024],prg00[3007:2992],prg00[2975:2960],prg00[2943:2928],prg00[2911:2896],prg00[2879:2864],prg00[2847:2832],
            prg00[2815:2800],prg00[2783:2768],prg00[2751:2736],prg00[2719:2704],prg00[2687:2672],prg00[2655:2640],prg00[2623:2608],prg00[2591:2576],
            prg00[2559:2544],prg00[2527:2512],prg00[2495:2480],prg00[2463:2448],prg00[2431:2416],prg00[2399:2384],prg00[2367:2352],prg00[2335:2320],
            prg00[2303:2288],prg00[2271:2256],prg00[2239:2224],prg00[2207:2192],prg00[2175:2160],prg00[2143:2128],prg00[2111:2096],prg00[2079:2064],
            prg00[2047:2032],prg00[2015:2000],prg00[1983:1968],prg00[1951:1936],prg00[1919:1904],prg00[1887:1872],prg00[1855:1840],prg00[1823:1808],
            prg00[1791:1776],prg00[1759:1744],prg00[1727:1712],prg00[1695:1680],prg00[1663:1648],prg00[1631:1616],prg00[1599:1584],prg00[1567:1552],
            prg00[1535:1520],prg00[1503:1488],prg00[1471:1456],prg00[1439:1424],prg00[1407:1392],prg00[1375:1360],prg00[1343:1328],prg00[1311:1296],
            prg00[1279:1264],prg00[1247:1232],prg00[1215:1200],prg00[1183:1168],prg00[1151:1136],prg00[1119:1104],prg00[1087:1072],prg00[1055:1040],
            prg00[1023:1008],prg00[ 991: 976],prg00[ 959: 944],prg00[ 927: 912],prg00[ 895: 880],prg00[ 863: 848],prg00[ 831: 816],prg00[ 799: 784],
            prg00[ 767: 752],prg00[ 735: 720],prg00[ 703: 688],prg00[ 671: 656],prg00[ 639: 624],prg00[ 607: 592],prg00[ 575: 560],prg00[ 543: 528],
            prg00[ 511: 496],prg00[ 479: 464],prg00[ 447: 432],prg00[ 415: 400],prg00[ 383: 368],prg00[ 351: 336],prg00[ 319: 304],prg00[ 287: 272],
            prg00[ 255: 240],prg00[ 223: 208],prg00[ 191: 176],prg00[ 159: 144],prg00[ 127: 112],prg00[  95:  80],prg00[  63:  48],prg00[  31:  16]};

   m_ebr_w16 #(.EBRADRWIDTH(EBRADRWIDTH),
               .prg0(pb0), .prg1(pb1), .prg2(pb2), .prg3(pb3), .prg4(pb4), .prg5(pb5), .prg6(pb6), .prg7(pb7) )
   ebrb 
     (/*AUTOINST*/
      // Outputs
      .DAT_O                            (eDAT_O[15:0]),
      // Inputs
      .B                                (B[15:0]),
      .Rai                              (Rai[EBRADRWIDTH-1:0]),
      .Wai                              (Wai[EBRADRWIDTH-1:0]),
      .clk                              (clk),
      .bmask                            (bmask[1:0]),
      .iwe                              (iwe));
   
   m_ebr_w16 #(.EBRADRWIDTH(EBRADRWIDTH),
               .prg0(ph0), .prg1(ph1), .prg2(ph2), .prg3(ph3), .prg4(ph4), .prg5(ph5), .prg6(ph6), .prg7(ph7) )
   ebrh
     (
      // Outputs
      .DAT_O                            (eDAT_O[31:16]),
      // Inputs
      .B                                (B[31:16]),
      .bmask                            (bmask[3:2]),
      /*AUTOINST*/
      // Inputs
      .Rai                              (Rai[EBRADRWIDTH-1:0]),
      .Wai                              (Wai[EBRADRWIDTH-1:0]),
      .clk                              (clk),
      .iwe                              (iwe));
   
endmodule
//MODE	DATA Width  Used WDATA/RDATA Bits
//0	16	    15, 14, 13, 12, 11, 10, 9, 8, 7, 6, 5, 4, 3, 2, 1, 0
//1	8	    14, 12, 10, 8, 6, 4, 2, 0
//2	4	    13, 9, 5, 1
//3	2	    11, 3

// Local Variables:
// verilog-library-directories:("."  )
// verilog-library-extensions:(".v" )
// End:
